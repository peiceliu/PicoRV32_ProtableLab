module back_fft_display(                                  //��ʾ�ַ���logo Ŀǰ������ӱ�������+���Σ������������ֿ��ܳ��ֵ��ӣ�����Ҫ��һ��ģ�鲢����Ҫ�ж����ȼ���
    input             lcd_pclk,     //ʱ��
    input             rst_n,        //��λ���͵�ƽ��Ч
                                    
    input      [10:0] pixel_xpos,   //���ص������
    input      [10:0] pixel_ypos,   //���ص������� 
    input      [1:0] wave_choose,
    output            wave_en   ,   //��ʾ��Щ�̶�������ʹ�� 
    output reg [23:0] pixel_data_wave,    //���ص�����,
    output            back_en   ,   //��ʾ��Щ�̶�������ʹ�� 
    output reg [23:0] pixel_data    //���ص�����,
);                                   
                                     
//parameter define                   
localparam PIC_X_START = 11'd10;     //ͼƬ��ʼ������� �Ϲ�ͬ����logo
localparam PIC_Y_START = 11'd10;     //ͼƬ��ʼ��������
localparam PIC_WIDTH   = 11'd64;    //ͼƬ���
localparam PIC_HEIGHT  = 11'd32;    //ͼƬ�߶�
       
localparam CHAR_X_START_bx= 11'd370;     //�ַ���ʼ������� ��ЯƵ���� 32x160
localparam CHAR_Y_START_bx= 11'd1;    //�ַ���ʼ��������
localparam CHAR_WIDTH_bx  = 11'd160;    //�ַ����, 48
localparam CHAR_HEIGHT = 11'd32;     //�ַ��߶�
wire  [10:0]  x_cnt_bx;       //�����������
wire  [10:0]  y_cnt_bx;       //�����������
assign  x_cnt_bx = pixel_xpos + 1'b1  - CHAR_X_START_bx; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_bx = pixel_ypos - CHAR_Y_START_bx; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_fdp= 11'd316;     //�ַ���ʼ������� ������ 96x32
localparam CHAR_Y_START_fdp= 11'd150;    //�ַ���ʼ��������
localparam CHAR_WIDTH_fdp  = 11'd96;    //�ַ����, 
wire  [10:0]  x_cnt_fdp;       //�����������
wire  [10:0]  y_cnt_fdp;       //�����������
assign  x_cnt_fdp = pixel_xpos + 1'b1  - CHAR_X_START_fdp; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_fdp = pixel_ypos - CHAR_Y_START_fdp; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_bxpl= 11'd10;     //�ַ���ʼ������� ����Ƶ�ʣ� 160x32
localparam CHAR_Y_START_bxpl= 11'd75;    //�ַ���ʼ��������
localparam CHAR_WIDTH_bxpl  = 11'd160;    //�ַ����, 
wire  [10:0]  x_cnt_bxpl;       //�����������
wire  [10:0]  y_cnt_bxpl;       //�����������
assign  x_cnt_bxpl = pixel_xpos + 1'b1  - CHAR_X_START_bxpl; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_bxpl = pixel_ypos - CHAR_Y_START_bxpl; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_bxzl= 11'd10;     //�ַ���ʼ������� �������ࣺ 160x32
localparam CHAR_Y_START_bxzl= 11'd43;    //�ַ���ʼ��������
localparam CHAR_WIDTH_bxzl  = 11'd160;    //�ַ����, 
wire  [10:0]  x_cnt_bxzl;       //�����������
wire  [10:0]  y_cnt_bxzl;       //�����������
assign  x_cnt_bxzl = pixel_xpos + 1'b1  - CHAR_X_START_bxzl; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_bxzl = pixel_ypos - CHAR_Y_START_bxzl; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_zxb= 11'd171;     //�ַ���ʼ������� ���Ҳ� 96x32
localparam CHAR_Y_START_zxb= 11'd43;    //�ַ���ʼ��������
localparam CHAR_WIDTH_zxb  = 11'd96;    //�ַ����, 
wire  [10:0]  x_cnt_zxb;       //�����������
wire  [10:0]  y_cnt_zxb;       //�����������
assign  x_cnt_zxb = pixel_xpos + 1'b1  - CHAR_X_START_zxb; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_zxb = pixel_ypos - CHAR_Y_START_zxb; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_jcb= 11'd171;     //�ַ���ʼ������� ��ݲ� 96x32
localparam CHAR_Y_START_jcb= 11'd43;    //�ַ���ʼ��������
localparam CHAR_WIDTH_jcb  = 11'd96;    //�ַ����, 
wire  [10:0]  x_cnt_jcb;       //�����������
wire  [10:0]  y_cnt_jcb;       //�����������
assign  x_cnt_jcb = pixel_xpos + 1'b1  - CHAR_X_START_jcb; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_jcb = pixel_ypos - CHAR_Y_START_jcb; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_sjb= 11'd171;     //�ַ���ʼ������� ���ǲ� 96x32
localparam CHAR_Y_START_sjb= 11'd43;    //�ַ���ʼ��������
localparam CHAR_WIDTH_sjb  = 11'd96;    //�ַ����, 
wire  [10:0]  x_cnt_sjb;       //�����������
wire  [10:0]  y_cnt_sjb;       //�����������
assign  x_cnt_sjb = pixel_xpos + 1'b1  - CHAR_X_START_sjb; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_sjb = pixel_ypos - CHAR_Y_START_sjb; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_fb= 11'd171;     //�ַ���ʼ������� ���� 96x32
localparam CHAR_Y_START_fb= 11'd43;    //�ַ���ʼ��������
localparam CHAR_WIDTH_fb  = 11'd96;    //�ַ����, 
wire  [10:0]  x_cnt_fb;       //�����������
wire  [10:0]  y_cnt_fb;       //�����������
assign  x_cnt_fb = pixel_xpos + 1'b1  - CHAR_X_START_fb; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_fb = pixel_ypos - CHAR_Y_START_fb; //���ص�������ַ�������ʼ�㴹ֱ����


localparam CHAR_X_START_FFT= 11'd350;     //�ַ���ʼ������� FFT:256   112x32
localparam CHAR_Y_START_FFT= 11'd43;    //�ַ���ʼ��������
localparam CHAR_WIDTH_FFT  = 11'd112;    //�ַ����, 
wire  [10:0]  x_cnt_FFT;       //�����������
wire  [10:0]  y_cnt_FFT;       //�����������
assign  x_cnt_FFT = pixel_xpos + 1'b1  - CHAR_X_START_FFT; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_FFT = pixel_ypos - CHAR_Y_START_FFT; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_ppbj= 11'd350;     //�ַ���ʼ������� Ƶ�ײ�����5   176x32
localparam CHAR_Y_START_ppbj= 11'd75;    //�ַ���ʼ��������
localparam CHAR_WIDTH_ppbj  = 11'd176;    //�ַ����, 
wire  [10:0]  x_cnt_ppbj;       //�����������
wire  [10:0]  y_cnt_ppbj;       //�����������
assign  x_cnt_ppbj = pixel_xpos + 1'b1  - CHAR_X_START_ppbj; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_ppbj = pixel_ypos - CHAR_Y_START_ppbj; //���ص�������ַ�������ʼ�㴹ֱ����


localparam CHAR_X_START_xsds= 11'd530;     //�ַ���ʼ������� ��ʾ������128   208x32
localparam CHAR_Y_START_xsds= 11'd43;    //�ַ���ʼ��������
localparam CHAR_WIDTH_xsds  = 11'd208;    //�ַ����, 
wire  [10:0]  x_cnt_xsds;       //�����������
wire  [10:0]  y_cnt_xsds;       //�����������
assign  x_cnt_xsds = pixel_xpos + 1'b1  - CHAR_X_START_xsds; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_xsds = pixel_ypos - CHAR_Y_START_xsds; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_sp= 11'd530;     //�ַ���ʼ������� ˮƽ��20/div   224x32
localparam CHAR_Y_START_sp= 11'd75;    //�ַ���ʼ��������
localparam CHAR_WIDTH_sp  = 11'd224;    //�ַ����, 
wire  [10:0]  x_cnt_sp;       //�����������
wire  [10:0]  y_cnt_sp;       //�����������
assign  x_cnt_sp = pixel_xpos + 1'b1  - CHAR_X_START_sp; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_sp = pixel_ypos - CHAR_Y_START_sp; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_0= 11'd47;     //�ַ���ʼ������� 0   16x32
localparam CHAR_Y_START_0= 11'd438;    //�ַ���ʼ��������
localparam CHAR_WIDTH_0  = 11'd16;    //�ַ����, 
wire  [10:0]  x_cnt_0;       //�����������
wire  [10:0]  y_cnt_0;       //�����������
assign  x_cnt_0 = pixel_xpos + 1'b1  - CHAR_X_START_0; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_0 = pixel_ypos - CHAR_Y_START_0; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_20= 11'd248;     //�ַ���ʼ������� 20   32x32
localparam CHAR_Y_START_20= 11'd438;    //�ַ���ʼ��������
localparam CHAR_WIDTH_20  = 11'd32;    //�ַ����, 
wire  [10:0]  x_cnt_20;       //�����������
wire  [10:0]  y_cnt_20;       //�����������
assign  x_cnt_20 = pixel_xpos + 1'b1  - CHAR_X_START_20; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_20 = pixel_ypos - CHAR_Y_START_20; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_40= 11'd448;     //�ַ���ʼ������� 40   32x32
localparam CHAR_Y_START_40= 11'd438;    //�ַ���ʼ��������
localparam CHAR_WIDTH_40  = 11'd32;    //�ַ����, 
wire  [10:0]  x_cnt_40;       //�����������
wire  [10:0]  y_cnt_40;       //�����������
assign  x_cnt_40 = pixel_xpos + 1'b1  - CHAR_X_START_40; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_40 = pixel_ypos - CHAR_Y_START_40; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_60= 11'd648;     //�ַ���ʼ������� 60/KHZ   96x32
localparam CHAR_Y_START_60= 11'd438;    //�ַ���ʼ��������
localparam CHAR_WIDTH_60  = 11'd96;    //�ַ����, 
wire  [10:0]  x_cnt_60;       //�����������
wire  [10:0]  y_cnt_60;       //�����������
assign  x_cnt_60 = pixel_xpos + 1'b1  - CHAR_X_START_60; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_60 = pixel_ypos - CHAR_Y_START_60; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_50= 11'd30;     //�ַ���ʼ������� 50   32x32
localparam CHAR_Y_START_50= 11'd370;    //�ַ���ʼ��������
localparam CHAR_WIDTH_50  = 11'd32;    //�ַ����, 
wire  [10:0]  x_cnt_50;       //�����������
wire  [10:0]  y_cnt_50;       //�����������
assign  x_cnt_50 = pixel_xpos + 1'b1  - CHAR_X_START_50; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_50 = pixel_ypos - CHAR_Y_START_50; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_100= 11'd14;     //�ַ���ʼ������� 100   48x32
localparam CHAR_Y_START_100= 11'd320;    //�ַ���ʼ��������
localparam CHAR_WIDTH_100  = 11'd48;    //�ַ����, 
wire  [10:0]  x_cnt_100;       //�����������
wire  [10:0]  y_cnt_100;       //�����������
assign  x_cnt_100 = pixel_xpos + 1'b1  - CHAR_X_START_100; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_100 = pixel_ypos - CHAR_Y_START_100; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_150= 11'd14;     //�ַ���ʼ������� 150   48x32
localparam CHAR_Y_START_150= 11'd270;    //�ַ���ʼ��������
localparam CHAR_WIDTH_150  = 11'd48;    //�ַ����, 
wire  [10:0]  x_cnt_150;       //�����������
wire  [10:0]  y_cnt_150;       //�����������
assign  x_cnt_150 = pixel_xpos + 1'b1  - CHAR_X_START_150; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_150 = pixel_ypos - CHAR_Y_START_150; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_200= 11'd14;     //�ַ���ʼ������� 200   48x32
localparam CHAR_Y_START_200= 11'd220;    //�ַ���ʼ��������
localparam CHAR_WIDTH_200  = 11'd48;    //�ַ����, 
wire  [10:0]  x_cnt_200;       //�����������
wire  [10:0]  y_cnt_200;       //�����������
assign  x_cnt_200 = pixel_xpos + 1'b1  - CHAR_X_START_200; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_200 = pixel_ypos - CHAR_Y_START_200; //���ص�������ַ�������ʼ�㴹ֱ����

localparam CHAR_X_START_256= 11'd64;     //�ַ���ʼ������� x256  64x32
localparam CHAR_Y_START_256= 11'd152;    //�ַ���ʼ��������
localparam CHAR_WIDTH_256  = 11'd64;    //�ַ����, 
wire  [10:0]  x_cnt_256;       //�����������
wire  [10:0]  y_cnt_256;       //�����������
assign  x_cnt_256 = pixel_xpos + 1'b1  - CHAR_X_START_256; //���ص�������ַ�������ʼ��ˮƽ����
assign  y_cnt_256 = pixel_ypos - CHAR_Y_START_256; //���ص�������ַ�������ʼ�㴹ֱ����


localparam BACK_COLOR  = 24'hffffff; //����ɫ����ɫ
//localparam CHAR_COLOR  = 24'hff0000; //�ַ���ɫ����ɫ
localparam BLUE   = 24'b00000000_00000000_11111111;     //RGB888 ��ɫ
localparam CHAR_COLOR  = 24'b00000000_00000000_00000000; //�ַ���ɫ����ɫ
//reg define
reg   [11:0]  rom_addr  ;  //ROM��ַ
wire          rom_rd_en ;  //ROM��ʹ���ź�
wire  [23:0]  rom_rd_data ;//ROM����
//*****************************************************
//**                    main code
//*****************************************************
assign  rom_rd_en = 1'b1;                  //��ʹ�����ߣ���һֱ��ROM����

reg [159:0] char_bx[31:0];
//��ЯƵ����
always @(posedge lcd_pclk) begin
    char_bx[0 ]  <=   160'h0000000000000000000000000000000000000000;
    char_bx[1 ]  <=   160'h0000000000000000000000000002010000000000;
    char_bx[2 ]  <=   160'h0080000001008000004000000001038000400000;
    char_bx[3 ]  <=   160'h00E000180180CC00006000080C01830000708000;
    char_bx[4 ]  <=   160'h00DFFFFC0100C6000061FFFC0600C20000E04000;
    char_bx[5 ]  <=   160'h0180180001018610006003000700843000C02000;
    char_bx[6 ]  <=   160'h018018000101FFF806600600031FFFF800C03000;
    char_bx[7 ]  <=   160'h0100182001030400066404000200C60001803840;
    char_bx[8 ]  <=   160'h030FFFF001230400067E04080010C62001801860;
    char_bx[9 ]  <=   160'h020C18303FF7042006607FFC0008C630030410E0;
    char_bx[10]  <=   160'h060C1830010FFFF006606018000CC670030400C0;
    char_bx[11]  <=   160'h070C1830010B0400066060180206C66003820080;
    char_bx[12]  <=   160'h0F0C183001130420066262187F06C6C007820180;
    char_bx[13]  <=   160'h0B0FFFF0010BFFF03FFF63980206C6800D820180;
    char_bx[14]  <=   160'h1B0C183001330400004063180200C70809810300;
    char_bx[15]  <=   160'h130C183001C3040000606318027FFFFC19810300;
    char_bx[16]  <=   160'h230C183003830418044063180200000011808600;
    char_bx[17]  <=   160'h430C18300F03FFFC06406318020000002180C600;
    char_bx[18]  <=   160'h030FFFF079030000064263180204004041804400;
    char_bx[19]  <=   160'h030C1830310200000C4763180207FFE001806C00;
    char_bx[20]  <=   160'h03001800010FFFC00C4663180206004001802800;
    char_bx[21]  <=   160'h0304100001004080184C6218021E004001803800;
    char_bx[22]  <=   160'h030210000100C188104C62180226004001803800;
    char_bx[23]  <=   160'h030130000100C3FC201807000266004001806C00;
    char_bx[24]  <=   160'h0300B000010081182030048002C7FFC001804600;
    char_bx[25]  <=   160'h0300E0000101801800600C600386004001808380;
    char_bx[26]  <=   160'h030070000103001800C0183807060040018301C0;
    char_bx[27]  <=   160'h0300DC00010600300180301C03060040018600F0;
    char_bx[28]  <=   160'h03030FC01F0C03300600600C0007FFC00188007E;
    char_bx[29]  <=   160'h030E03FC073001E0080180040006004001B00030;
    char_bx[30]  <=   160'h02F00038024000C0300600040006004001400000;
    char_bx[31]  <=   160'h0000000000000000000000000000000000000000;
    end 
 reg [223:0] char_sp[31:0];
    //ˮƽ��20/div
always @(posedge lcd_pclk) begin
        char_sp[0 ]  <=   224'h00000000000000000000000000000000000000000000000000000000;
        char_sp[1 ]  <=   224'h00000000000000000000000000000000000000000000000000000000;
        char_sp[2 ]  <=   224'h00038000000000000000000000000000000100000000000000000000;
        char_sp[3 ]  <=   224'h0003E000000000600000000000000000000180000002000000000000;
        char_sp[4 ]  <=   224'h000380000FFFFFF00000000000000000000180000006000000000000;
        char_sp[5 ]  <=   224'h00038000000180000000000000000000000180000004000800000000;
        char_sp[6 ]  <=   224'h0003C000000180000000000007E003C000018060000C007801800000;
        char_sp[7 ]  <=   224'h0003C0600201818000000000083806200001FFF00008001803C00000;
        char_sp[8 ]  <=   224'h0003C0F0010181C00000000010180C30000180000018001801800000;
        char_sp[9 ]  <=   224'h0003C1F000C1818000000000200C1818000180000010001800000000;
        char_sp[10]  <=   224'h003BC3E000C1830000000000200C1818000180000030001800000000;
        char_sp[11]  <=   224'h3FFFE78000E1820000000000300C1808000180000020001800000000;
        char_sp[12]  <=   224'h187BEF000061840000000000300C300C010180800060001800800000;
        char_sp[13]  <=   224'h007BFC000061880000000000000C300C01FFFFC0004007D81F807C3E;
        char_sp[14]  <=   224'h0073F80000218800000000000018300C0180018000C00C380180180C;
        char_sp[15]  <=   224'h00F3F80000019018000000000018300C018001800080181801801808;
        char_sp[16]  <=   224'h00F3F8007FFFFFFC000000000030300C018001800180181801801818;
        char_sp[17]  <=   224'h00E3DC0000018000070000000060300C018001800100301801800C10;
        char_sp[18]  <=   224'h01E3DE00000180000F00000000C0300C018001800300301801800C10;
        char_sp[19]  <=   224'h01C3CE00000180000F0000000180300C018001800200301801800420;
        char_sp[20]  <=   224'h03C3CF0000018000070000000300300C01FFFF800600301801800620;
        char_sp[21]  <=   224'h0383C78000018000000000000200300C018001800400301801800620;
        char_sp[22]  <=   224'h0703C3C0000180000000000004041808018001000C00301801800340;
        char_sp[23]  <=   224'h0703C3E0000180000000000008041818000000000800301801800340;
        char_sp[24]  <=   224'h0E03C1F80001800000000000100418180010204018001018018003C0;
        char_sp[25]  <=   224'h1C03C0FE0001800007000000200C0C30020830601000183801800180;
        char_sp[26]  <=   224'h3803C07E000180000F0000003FF80620020C183030000C5E01800180;
        char_sp[27]  <=   224'h7023C038000180000F0000003FF803C0060C1838200007901FF80100;
        char_sp[28]  <=   224'h607F80000001800006000000000000000C0618186000000000000000;
        char_sp[29]  <=   224'h000F80000001800000000000000000001C0408184000000000000000;
        char_sp[30]  <=   224'h00070000000100000000000000000000180400100000000000000000;
        char_sp[31]  <=   224'h00000000000000000000000000000000000000000000000000000000;
        end 

reg [95:0] char_fdp[31:0];
 //������
always @(posedge lcd_pclk) begin
        char_fdp[0 ]  <=   96'h000000000000000000000000;
        char_fdp[1 ]  <=   96'h000000000000000000020100;
        char_fdp[2 ]  <=   96'h038000000001000000010380;
        char_fdp[3 ]  <=   96'h03C0001C0000C0000C018300;
        char_fdp[4 ]  <=   96'h038FFFFE0000E0100600C200;
        char_fdp[5 ]  <=   96'h038600000400403807008430;
        char_fdp[6 ]  <=   96'h0380000007FFFFFC031FFFF8;
        char_fdp[7 ]  <=   96'h3398C060060404000200C600;
        char_fdp[8 ]  <=   96'h3FFCFFF0060707000010C620;
        char_fdp[9 ]  <=   96'h3BB8E0F0060606000008C630;
        char_fdp[10]  <=   96'h3BB8E0E006060630000CC670;
        char_fdp[11]  <=   96'h3BB8E0E007FFFFF80206C660;
        char_fdp[12]  <=   96'h3BB8E0E0060606007F06C6C0;
        char_fdp[13]  <=   96'h3BB8FFE0060606000206C680;
        char_fdp[14]  <=   96'h3BB8E0E0060606000200C708;
        char_fdp[15]  <=   96'h3BB8E0C006060600027FFFFC;
        char_fdp[16]  <=   96'h3BBB00180607FE0002000000;
        char_fdp[17]  <=   96'h3BBBFFFC0606060002000000;
        char_fdp[18]  <=   96'h3BBB8E3C0400010002040040;
        char_fdp[19]  <=   96'h3BBB8E3C043FFF800207FFE0;
        char_fdp[20]  <=   96'h3BBB8E3C0C04038002060040;
        char_fdp[21]  <=   96'h3BFB8E3C0C020700021E0040;
        char_fdp[22]  <=   96'h3BFBFFFC0C03060002260040;
        char_fdp[23]  <=   96'h3BB38E3C08010C0002660040;
        char_fdp[24]  <=   96'h33838E3C0800D80002C7FFC0;
        char_fdp[25]  <=   96'h03838E3C1800700003860040;
        char_fdp[26]  <=   96'h03838E3C1000F80007060040;
        char_fdp[27]  <=   96'h03838E3C10039E0003060040;
        char_fdp[28]  <=   96'h0383FFFC200E07F80007FFC0;
        char_fdp[29]  <=   96'h0383803C207000F800060040;
        char_fdp[30]  <=   96'h038380384780001000060040;
        char_fdp[31]  <=   96'h038300100000000000000000;
        end 
reg [159:0] char_bxzl[31:0];
//�������ࣺ
always @(posedge lcd_pclk) begin
    char_bxzl[0 ]  <=   160'h0000000000000000000000000000000000000000;
    char_bxzl[1 ]  <=   160'h0000000000000000000000000000000000000000;
    char_bxzl[2 ]  <=   160'h00001C0000000000000004000001800000000000;
    char_bxzl[3 ]  <=   160'h0E001C0000000020001807000101C18000000000;
    char_bxzl[4 ]  <=   160'h0F001C0000006070007C060000C181C000000000;
    char_bxzl[5 ]  <=   160'h07801C001FFFF0E00FC006000071830000000000;
    char_bxzl[6 ]  <=   160'h03801C00018200C030C006000031860000000000;
    char_bxzl[7 ]  <=   160'h039C1C380182018000C006000031840000000000;
    char_bxzl[8 ]  <=   160'h003FFFFC0182030000C006000021881800000000;
    char_bxzl[9 ]  <=   160'h003E1C7C0182060000C106103FFFFFFC00000000;
    char_bxzl[10]  <=   160'h707E1C700182040000C9FFF80007800000000000;
    char_bxzl[11]  <=   160'h3C7E1CE0018208003FFF8618000DF00000000000;
    char_bxzl[12]  <=   160'h1CFE1CC00182101000C1861800198E0000000000;
    char_bxzl[13]  <=   160'h1EDE1C000182603801C18618003183C000000000;
    char_bxzl[14]  <=   160'h0EDE1C603FFFF07001C18618006180F000000000;
    char_bxzl[15]  <=   160'h0DDFFFF0018200C001E1861801C1807000000000;
    char_bxzl[16]  <=   160'h019EC0F00182018003D986180301003000000000;
    char_bxzl[17]  <=   160'h039EC0E00182030002DD86181C03001007000000;
    char_bxzl[18]  <=   160'h039CE1E00182060006CDFFF8200380080F000000;
    char_bxzl[19]  <=   160'h071C61C00182080004C18618000300180F000000;
    char_bxzl[20]  <=   160'h071C7380010230080CC186107FFFFFFC07000000;
    char_bxzl[21]  <=   160'h7E1C37800302001C18C006000002400000000000;
    char_bxzl[22]  <=   160'h7E1C3F000302003810C006000006200000000000;
    char_bxzl[23]  <=   160'h1E381E000202007020C006000006300000000000;
    char_bxzl[24]  <=   160'h0E381E00060200C040C00600000C180000000000;
    char_bxzl[25]  <=   160'h1E703F800402018000C0060000180C0007000000;
    char_bxzl[26]  <=   160'h1E70F7C00C02030000C00600003807000F000000;
    char_bxzl[27]  <=   160'h1EE1E3F008020E0000C00600007003E00F000000;
    char_bxzl[28]  <=   160'h1FC7C0FE1002180000C0060001C000FE06000000;
    char_bxzl[29]  <=   160'h1F9F007C2004600000C006000700007000000000;
    char_bxzl[30]  <=   160'h0378001000008000008004003800000000000000;
    char_bxzl[31]  <=   160'h0000000000000000000000000000000000000000;
    end 
reg [159:0] char_bxpl[31:0];
    //����Ƶ�ʣ�
always @(posedge lcd_pclk) begin
        char_bxpl[0 ]  <=   160'h0000000000000000000000000000000000000000;
        char_bxpl[1 ]  <=   160'h0000000000000000000000000000000000000000;
        char_bxpl[2 ]  <=   160'h00001C0000000000004000000002000000000000;
        char_bxpl[3 ]  <=   160'h0E001C0000000020006000080003800000000000;
        char_bxpl[4 ]  <=   160'h0F001C00000060700061FFFC0001800000000000;
        char_bxpl[5 ]  <=   160'h07801C001FFFF0E0006003000001802000000000;
        char_bxpl[6 ]  <=   160'h03801C00018200C0066006001FFFFFF000000000;
        char_bxpl[7 ]  <=   160'h039C1C3801820180066404000003000000000000;
        char_bxpl[8 ]  <=   160'h003FFFFC01820300067E04080003000000000000;
        char_bxpl[9 ]  <=   160'h003E1C7C0182060006607FFC0C06104000000000;
        char_bxpl[10]  <=   160'h707E1C700182040006606018070C38E000000000;
        char_bxpl[11]  <=   160'h3C7E1CE001820800066060180398318000000000;
        char_bxpl[12]  <=   160'h1CFE1CC00182101006626218013FE30000000000;
        char_bxpl[13]  <=   160'h1EDE1C00018260383FFF63980138C40000000000;
        char_bxpl[14]  <=   160'h0EDE1C603FFFF070004063180001800000000000;
        char_bxpl[15]  <=   160'h0DDFFFF0018200C0006063180043020000000000;
        char_bxpl[16]  <=   160'h019EC0F00182018004406318008621C000000000;
        char_bxpl[17]  <=   160'h039EC0E00182030006406318030818E007000000;
        char_bxpl[18]  <=   160'h039CE1E001820600064263180E3FFC300F000000;
        char_bxpl[19]  <=   160'h071C61C0018208000C4763181C3D0C300F000000;
        char_bxpl[20]  <=   160'h071C7380010230080C4663180801880007000000;
        char_bxpl[21]  <=   160'h7E1C37800302001C184C62180001800000000000;
        char_bxpl[22]  <=   160'h7E1C3F0003020038104C62180001801800000000;
        char_bxpl[23]  <=   160'h1E381E0002020070201807003FFFFFFC00000000;
        char_bxpl[24]  <=   160'h0E381E00060200C0203004800001800000000000;
        char_bxpl[25]  <=   160'h1E703F800402018000600C600001800007000000;
        char_bxpl[26]  <=   160'h1E70F7C00C02030000C01838000180000F000000;
        char_bxpl[27]  <=   160'h1EE1E3F008020E000180301C000180000F000000;
        char_bxpl[28]  <=   160'h1FC7C0FE100218000600600C0001800006000000;
        char_bxpl[29]  <=   160'h1F9F007C20046000080180040001800000000000;
        char_bxpl[30]  <=   160'h0378001000008000300600040001000000000000;
        char_bxpl[31]  <=   160'h0000000000000000000000000000000000000000;
        end 
reg [95:0] char_zxb[31:0];
//���Ҳ�
always @(posedge lcd_pclk) begin
            char_zxb[0 ]  <=   96'h000000000000000000000000;
            char_zxb[1 ]  <=   96'h000000000000000000000000;
            char_zxb[2 ]  <=   96'h000000000000200000001800;
            char_zxb[3 ]  <=   96'h00000030002018000C001800;
            char_zxb[4 ]  <=   96'h000000781FF00C0006001800;
            char_zxb[5 ]  <=   96'h0FFFFFFC00200C0003001800;
            char_zxb[6 ]  <=   96'h0601E00000200C1803001800;
            char_zxb[7 ]  <=   96'h0001E0000027FFFC01081810;
            char_zxb[8 ]  <=   96'h0001E00000200800001FFFF8;
            char_zxb[9 ]  <=   96'h0001E00000201C00002C1838;
            char_zxb[10]  <=   96'h0001E00000201800202C1820;
            char_zxb[11]  <=   96'h0001E0000FE03000184C1840;
            char_zxb[12]  <=   96'h01E1E000082020401C4C1800;
            char_zxb[13]  <=   96'h01F1E040080060E00C4C1800;
            char_zxb[14]  <=   96'h01E1E0E0080040C00C8C1820;
            char_zxb[15]  <=   96'h01E1FFF018008180008FFFF0;
            char_zxb[16]  <=   96'h01E1E00018011F00010C8060;
            char_zxb[17]  <=   96'h01E1E0001821E300010C80C0;
            char_zxb[18]  <=   96'h01E1E0003FF10600010C40C0;
            char_zxb[19]  <=   96'h01E1E00010200C00020C4180;
            char_zxb[20]  <=   96'h01E1E0000020080002082180;
            char_zxb[21]  <=   96'h01E1E0000060180006083300;
            char_zxb[22]  <=   96'h01E1E000006030C03C181E00;
            char_zxb[23]  <=   96'h01E1E000006060600C100E00;
            char_zxb[24]  <=   96'h01E1E0000060C0300C100C00;
            char_zxb[25]  <=   96'h01E1E000006180380C201F00;
            char_zxb[26]  <=   96'h01E1E0300063FFD80C607380;
            char_zxb[27]  <=   96'h01E1E07800C3F0180C40C1E0;
            char_zxb[28]  <=   96'h7FFFFFFC1FC100080C83807C;
            char_zxb[29]  <=   96'h3000000003800000050E0038;
            char_zxb[30]  <=   96'h000000000300000002300000;
            char_zxb[31]  <=   96'h000000000000000000000000;
            end 
 reg [95:0] char_jcb[31:0];
//��ݲ�
 always @(posedge lcd_pclk) begin
 char_jcb[0 ]  <=   96'h000000000000000000000000;
 char_jcb[1 ]  <=   96'h000000000000000000000000;
 char_jcb[2 ]  <=   96'h038000100000800000001800;
 char_jcb[3 ]  <=   96'h07C3003C0000C0000C001800;
 char_jcb[4 ]  <=   96'h0783FFFC0180C00006001800;
 char_jcb[5 ]  <=   96'h0703803801C0C00003001800;
 char_jcb[6 ]  <=   96'h073B80380180C0C003001800;
 char_jcb[7 ]  <=   96'h0FFF80380180FFE001081810;
 char_jcb[8 ]  <=   96'h0E0380380180C000001FFFF8;
 char_jcb[9 ]  <=   96'h0E03FFF80180C000002C1838;
 char_jcb[10]  <=   96'h1C0380380180C000202C1820;
 char_jcb[11]  <=   96'h183B87800180C018184C1840;
 char_jcb[12]  <=   96'h3FFB87003FFFFFFC1C4C1800;
 char_jcb[13]  <=   96'h33838700000100000C4C1800;
 char_jcb[14]  <=   96'h6383871C0001C0000C8C1820;
 char_jcb[15]  <=   96'h6383FFFE0201C040008FFFF0;
 char_jcb[16]  <=   96'h0383870003018070010C8060;
 char_jcb[17]  <=   96'h039B870003018060010C80C0;
 char_jcb[18]  <=   96'h7FFF870003038060010C40C0;
 char_jcb[19]  <=   96'h3383C73803034060020C4180;
 char_jcb[20]  <=   96'h0383FFFC0302206002082180;
 char_jcb[21]  <=   96'h0387E0380306186006083300;
 char_jcb[22]  <=   96'h0387E038030C1C603C181E00;
 char_jcb[23]  <=   96'h03BFE03803080C600C100E00;
 char_jcb[24]  <=   96'h03FEE038031006600C100C00;
 char_jcb[25]  <=   96'h03EEE038036004600C201F00;
 char_jcb[26]  <=   96'h03DCE038038000600C607380;
 char_jcb[27]  <=   96'h039CE038030000600C40C1E0;
 char_jcb[28]  <=   96'h0338FFF807FFFFE00C83807C;
 char_jcb[29]  <=   96'h0070E03802000060050E0038;
 char_jcb[30]  <=   96'h0060E0200000004002300000;
 char_jcb[31]  <=   96'h000000000000000000000000;
 end 
 reg [95:0] char_sjb[31:0];
 //���ǲ�
  always @(posedge lcd_pclk) begin
  char_sjb[0 ]  <=   96'h000000000000000000000000;
  char_sjb[1 ]  <=   96'h000000000000000000000000;
  char_sjb[2 ]  <=   96'h000000000010000000001800;
  char_sjb[3 ]  <=   96'h00000000001C00000C001800;
  char_sjb[4 ]  <=   96'h000000000018000006001800;
  char_sjb[5 ]  <=   96'h000000600030080003001800;
  char_sjb[6 ]  <=   96'h000000F0007FFC0003001800;
  char_sjb[7 ]  <=   96'h1FFFFFF80060180001081810;
  char_sjb[8 ]  <=   96'h0C00000000C03000001FFFF8;
  char_sjb[9 ]  <=   96'h0000000001802060002C1838;
  char_sjb[10]  <=   96'h0000000001FFFFF0202C1820;
  char_sjb[11]  <=   96'h0000000003C0C060184C1840;
  char_sjb[12]  <=   96'h0000000004C0C0601C4C1800;
  char_sjb[13]  <=   96'h0000000008C0C0600C4C1800;
  char_sjb[14]  <=   96'h0000018030C0C0600C8C1820;
  char_sjb[15]  <=   96'h000003C000FFFFE0008FFFF0;
  char_sjb[16]  <=   96'h07FFFFE000C0C060010C8060;
  char_sjb[17]  <=   96'h0300000000C0C060010C80C0;
  char_sjb[18]  <=   96'h0000000000C0C060010C40C0;
  char_sjb[19]  <=   96'h0000000000C0C060020C4180;
  char_sjb[20]  <=   96'h0000000000FFFFE002082180;
  char_sjb[21]  <=   96'h000000000080C06006083300;
  char_sjb[22]  <=   96'h000000000080C0603C181E00;
  char_sjb[23]  <=   96'h000000000180C0600C100E00;
  char_sjb[24]  <=   96'h000000000180C0600C100C00;
  char_sjb[25]  <=   96'h000000180300C0600C201F00;
  char_sjb[26]  <=   96'h0000003C0200C0600C607380;
  char_sjb[27]  <=   96'h7FFFFFFE0600C0600C40C1E0;
  char_sjb[28]  <=   96'h300000000C00C7E00C83807C;
  char_sjb[29]  <=   96'h00000000100081E0050E0038;
  char_sjb[30]  <=   96'h000000002000008002300000;
  char_sjb[31]  <=   96'h000000000000000000000000;
  end 
  reg [95:0] char_fb[31:0];
// ����
always @(posedge lcd_pclk) begin
    char_fb[0 ]  <=   96'h000000000000000000000000;
    char_fb[1 ]  <=   96'h000000000000000000000000;
    char_fb[2 ]  <=   96'h000000060000000018000000;
    char_fb[3 ]  <=   96'h0000000380000C0018000000;
    char_fb[4 ]  <=   96'h000000018000060018000000;
    char_fb[5 ]  <=   96'h00000001C000030018000000;
    char_fb[6 ]  <=   96'h000000008000030018000000;
    char_fb[7 ]  <=   96'h000000000018010818100000;
    char_fb[8 ]  <=   96'h00003FFFFFFC001FFFF80000;
    char_fb[9 ]  <=   96'h000000060000002C18380000;
    char_fb[10]  <=   96'h000000060000202C18200000;
    char_fb[11]  <=   96'h000000060000184C18400000;
    char_fb[12]  <=   96'h0000000600001C4C18000000;
    char_fb[13]  <=   96'h0000000600800C4C18000000;
    char_fb[14]  <=   96'h00000007FFC00C8C18200000;
    char_fb[15]  <=   96'h000000060180008FFFF00000;
    char_fb[16]  <=   96'h000000040180010C80600000;
    char_fb[17]  <=   96'h0000000C0180010C80C00000;
    char_fb[18]  <=   96'h0000000C0180010C40C00000;
    char_fb[19]  <=   96'h000000080300020C41800000;
    char_fb[20]  <=   96'h000000180300020821800000;
    char_fb[21]  <=   96'h000000100300060833000000;
    char_fb[22]  <=   96'h0000003003003C181E000000;
    char_fb[23]  <=   96'h0000002003000C100E000000;
    char_fb[24]  <=   96'h0000006003000C100C000000;
    char_fb[25]  <=   96'h000000C002000C201F000000;
    char_fb[26]  <=   96'h0000018006000C6073800000;
    char_fb[27]  <=   96'h0000030186000C40C1E00000;
    char_fb[28]  <=   96'h000004007E000C83807C0000;
    char_fb[29]  <=   96'h000018003C00050E00380000;
    char_fb[30]  <=   96'h000020003000023000000000;
    char_fb[31]  <=   96'h000000000000000000000000;
    end 
    reg [175:0] char_ppbj[31:0];  
 //Ƶ�ײ�����5
always @(posedge lcd_pclk) begin
        char_ppbj[0 ]  <=   176'h00000000000000000000000000000000000000000000;
        char_ppbj[1 ]  <=   176'h00000000000201000000000000000000000000000000;
        char_ppbj[2 ]  <=   176'h00E00008000103800000800000010200000000000000;
        char_ppbj[3 ]  <=   176'h00F0001C0C0183000000C0000401C380000000000000;
        char_ppbj[4 ]  <=   176'h00E3FFFE0600C2000000800006018300000000000000;
        char_ppbj[5 ]  <=   176'h0CE18700070084300180800003018300000000000000;
        char_ppbj[6 ]  <=   176'h0FE00700031FFFF801C0804001818300000000000FFC;
        char_ppbj[7 ]  <=   176'h0EEE06000200C6000180FFE001018330000000000FFC;
        char_ppbj[8 ]  <=   176'h0EFFCE1C0010C62001808000003FFFF8000000001000;
        char_ppbj[9 ]  <=   176'h0EE0FFFE0008C6300180800000018300000000001000;
        char_ppbj[10]  <=   176'h0EE0E01C000CC6700180800000018300000000001000;
        char_ppbj[11]  <=   176'h0EE0E01C0206C6600180800000018300000000001000;
        char_ppbj[12]  <=   176'h0EE7E71C7F06C6C00180801801018300000000001000;
        char_ppbj[13]  <=   176'h7FFFE7DC0206C6803FFFFFFC7F818300000000001000;
        char_ppbj[14]  <=   176'h30E0E79C0200C70800010000030183000000000013E0;
        char_ppbj[15]  <=   176'h00F0E79C027FFFFC0000C00003018318000000001430;
        char_ppbj[16]  <=   176'h06E0E79C0200000000008000033FFFFC000000001818;
        char_ppbj[17]  <=   176'h0FE0E79C020000000040806003018300070000001008;
        char_ppbj[18]  <=   176'h0FE7E79C0204004000F08070030183000F000000000C;
        char_ppbj[19]  <=   176'h0EE7E71C0207FFE000C080E0030183000F000000000C;
        char_ppbj[20]  <=   176'h1CEFE71C02060040018081C00301030007000000000C;
        char_ppbj[21]  <=   176'h1CFEE71C021E0040030083000303030000000000000C;
        char_ppbj[22]  <=   176'h38FCE71C02260040020086000302030000000000300C;
        char_ppbj[23]  <=   176'h303CCF90026600400400DC000304030000000000300C;
        char_ppbj[24]  <=   176'h60780FE002C7FFC00801380003080300000000002018;
        char_ppbj[25]  <=   176'h00F01EF0038600401000E00004900300070000002018;
        char_ppbj[26]  <=   176'h01E03C7C070600400001C000186002000F0000001830;
        char_ppbj[27]  <=   176'h03C0783E0306004000070000303800020F00000007C0;
        char_ppbj[28]  <=   176'h0F00F01E0007FFC000380000300FFFFC060000000000;
        char_ppbj[29]  <=   176'h1E03C00E0006004003C000000001FFF0000000000000;
        char_ppbj[30]  <=   176'h700F000C000600403C00000000000000000000000000;
        char_ppbj[31]  <=   176'h00000000000000000000000000000000000000000000;
        end 
 reg [111:0] char_FFT[31:0];  
//FFT:256
always @(posedge lcd_pclk) begin
char_FFT[0 ]  <=   112'h0000000000000000000000000000;
char_FFT[1 ]  <=   112'h0000000000000000000000000000;
char_FFT[2 ]  <=   112'h0000000000000000000000000000;
char_FFT[3 ]  <=   112'h0000000000000000000000000000;
char_FFT[4 ]  <=   112'h0000000000000000000000000000;
char_FFT[5 ]  <=   112'h0000000000000000000000000000;
char_FFT[6 ]  <=   112'hFFFE7FFC3FFC000007E00FFC01E0;
char_FFT[7 ]  <=   112'h3C3E181C3184000008380FFC0618;
char_FFT[8 ]  <=   112'h3C0E180421860000101810000C18;
char_FFT[9 ]  <=   112'h3C07180241820000200C10000818;
char_FFT[10]  <=   112'h3C03180241820000200C10001800;
char_FFT[11]  <=   112'h3C00180001800000300C10001000;
char_FFT[12]  <=   112'h3C00180001800000300C10001000;
char_FFT[13]  <=   112'h3C38181001800180000C10003000;
char_FFT[14]  <=   112'h3C381810018003C0001813E033E0;
char_FFT[15]  <=   112'h3C381830018003C0001814303630;
char_FFT[16]  <=   112'h3FF81FF001800180003018183818;
char_FFT[17]  <=   112'h3C78183001800000006010083808;
char_FFT[18]  <=   112'h3C3818100180000000C0000C300C;
char_FFT[19]  <=   112'h3C381810018000000180000C300C;
char_FFT[20]  <=   112'h3C381810018000000300000C300C;
char_FFT[21]  <=   112'h3C001800018000000200000C300C;
char_FFT[22]  <=   112'h3C001800018000000404300C300C;
char_FFT[23]  <=   112'h3C001800018000000804300C180C;
char_FFT[24]  <=   112'h3C00180001800180100420181808;
char_FFT[25]  <=   112'h3C001800018003C0200C20180C18;
char_FFT[26]  <=   112'h3C001800018003C03FF818300E30;
char_FFT[27]  <=   112'hFF007E0007E001803FF807C003E0;
char_FFT[28]  <=   112'h0000000000000000000000000000;
char_FFT[29]  <=   112'h0000000000000000000000000000;
char_FFT[30]  <=   112'h0000000000000000000000000000;
char_FFT[31]  <=   112'h0000000000000000000000000000;
end 
reg [207:0] char_xsds[31:0];  
//��ʾ������128
always @(posedge lcd_pclk) begin
char_xsds[0 ]  <=   208'h0000000000000000000000000000000000000000000000000000;
char_xsds[1 ]  <=   208'h0000000000000000000000000000000000000000000000000000;
char_xsds[2 ]  <=   208'h0000000000000000000100000060080000000000000000000000;
char_xsds[3 ]  <=   208'h01800380000000800001800000700E0000000000000000000000;
char_xsds[4 ]  <=   208'h01FFFFC0000000C0000180000C618C0000000000000000000000;
char_xsds[5 ]  <=   208'h01C0038003FFFFE0000180000663180000000000000000000000;
char_xsds[6 ]  <=   208'h01C0038000000000000180600766180000000000008007E007E0;
char_xsds[7 ]  <=   208'h01C00380000000000001FFF00264100000000000018008380C30;
char_xsds[8 ]  <=   208'h01C00380000000000001800000691008000000001F8010181818;
char_xsds[9 ]  <=   208'h01FFFF8000000000000180003FFFFFFC000000000180200C300C;
char_xsds[10]  <=   208'h01C00380000000000001800000E03060000000000180200C300C;
char_xsds[11]  <=   208'h01C00380000000000001800001F83060000000000180300C300C;
char_xsds[12]  <=   208'h01C003800000001801018080016E7060000000000180300C380C;
char_xsds[13]  <=   208'h01C003803FFFFFFC01FFFFC002665060000000000180000C3808;
char_xsds[14]  <=   208'h01FFFF8000018000018001800462904000000000018000181E18;
char_xsds[15]  <=   208'h01C0038000018000018001801860904000000000018000180F20;
char_xsds[16]  <=   208'h019863000001800001800180204108C0000000000180003007C0;
char_xsds[17]  <=   208'h001E7860006188000180018000E008C0070000000180006018F0;
char_xsds[18]  <=   208'h181E787000F184000180018000C208C00F000000018000C03078;
char_xsds[19]  <=   208'h1C1C78F800C18300018001803FFF0C800F000000018001803038;
char_xsds[20]  <=   208'h0F1C78F001C1818001FFFF8001860D800700000001800300601C;
char_xsds[21]  <=   208'h079C79E0018180C001800180010605800000000001800200600C;
char_xsds[22]  <=   208'h07DC7BC0030180E001800100030C07000000000001800404600C;
char_xsds[23]  <=   208'h03DC7B800601807000000000038C07000000000001800804600C;
char_xsds[24]  <=   208'h03DC7F000C01803800102040007807000000000001801004600C;
char_xsds[25]  <=   208'h01DC7E000801801802083060003F0D80070000000180200C3018;
char_xsds[26]  <=   208'h001C7C3010018010020C183000E318E00F00000003C03FF81830;
char_xsds[27]  <=   208'h001C787820618000060C1838018130700F0000001FF83FF807C0;
char_xsds[28]  <=   208'h7FFFFFFC001F80000C0618180600C03E06000000000000000000;
char_xsds[29]  <=   208'h38000000000700001C0408183801001000000000000000000000;
char_xsds[30]  <=   208'h0000000000020000180400100006000000000000000000000000;
char_xsds[31]  <=   208'h0000000000000000000000000000000000000000000000000000;
end 
reg [15:0] char_0[31:0]; 
//0
always @(posedge lcd_pclk) begin
    char_0[0 ]  <=   16'h0000;
    char_0[1 ]  <=   16'h0000;
    char_0[2 ]  <=   16'h0000;
    char_0[3 ]  <=   16'h0000;
    char_0[4 ]  <=   16'h0000;
    char_0[5 ]  <=   16'h0000;
    char_0[6 ]  <=   16'h07E0;
    char_0[7 ]  <=   16'h0FF0;
    char_0[8 ]  <=   16'h1C38;
    char_0[9 ]  <=   16'h3C3C;
    char_0[10]  <=   16'h3C1C;
    char_0[11]  <=   16'h781C;
    char_0[12]  <=   16'h781E;
    char_0[13]  <=   16'h781E;
    char_0[14]  <=   16'h781E;
    char_0[15]  <=   16'h781E;
    char_0[16]  <=   16'h781E;
    char_0[17]  <=   16'h781E;
    char_0[18]  <=   16'h781E;
    char_0[19]  <=   16'h781E;
    char_0[20]  <=   16'h781E;
    char_0[21]  <=   16'h781E;
    char_0[22]  <=   16'h781C;
    char_0[23]  <=   16'h383C;
    char_0[24]  <=   16'h3C3C;
    char_0[25]  <=   16'h1C38;
    char_0[26]  <=   16'h0FF0;
    char_0[27]  <=   16'h07E0;
    char_0[28]  <=   16'h0000;
    char_0[29]  <=   16'h0000;
    char_0[30]  <=   16'h0000;
    char_0[31]  <=   16'h0000;
end 
reg [31:0] char_50[31:0]; 
//50
always @(posedge lcd_pclk) begin
    char_50[0 ]  <=   32'h00000000;
    char_50[1 ]  <=   32'h00000000;
    char_50[2 ]  <=   32'h00000000;
    char_50[3 ]  <=   32'h00000000;
    char_50[4 ]  <=   32'h00000000;
    char_50[5 ]  <=   32'h00000000;
    char_50[6 ]  <=   32'h1FFC03C0;
    char_50[7 ]  <=   32'h1FFC0620;
    char_50[8 ]  <=   32'h38000C30;
    char_50[9 ]  <=   32'h38001818;
    char_50[10]  <=   32'h38001818;
    char_50[11]  <=   32'h38001808;
    char_50[12]  <=   32'h3800300C;
    char_50[13]  <=   32'h39C0300C;
    char_50[14]  <=   32'h3FF0300C;
    char_50[15]  <=   32'h3E78300C;
    char_50[16]  <=   32'h383C300C;
    char_50[17]  <=   32'h381C300C;
    char_50[18]  <=   32'h001E300C;
    char_50[19]  <=   32'h001E300C;
    char_50[20]  <=   32'h001E300C;
    char_50[21]  <=   32'h381E300C;
    char_50[22]  <=   32'h781E1808;
    char_50[23]  <=   32'h781C1818;
    char_50[24]  <=   32'h781C1818;
    char_50[25]  <=   32'h383C0C30;
    char_50[26]  <=   32'h1E780620;
    char_50[27]  <=   32'h0FF003C0;
    char_50[28]  <=   32'h00000000;
    char_50[29]  <=   32'h00000000;
    char_50[30]  <=   32'h00000000;
    char_50[31]  <=   32'h00000000;
end 
reg [31:0] char_20[31:0]; 
//20
always @(posedge lcd_pclk) begin
    char_20[0 ]  <=   32'h00000000;
    char_20[1 ]  <=   32'h00000000;
    char_20[2 ]  <=   32'h00000000;
    char_20[3 ]  <=   32'h00000000;
    char_20[4 ]  <=   32'h00000000;
    char_20[5 ]  <=   32'h00000000;
    char_20[6 ]  <=   32'h0FF003C0;
    char_20[7 ]  <=   32'h1E780620;
    char_20[8 ]  <=   32'h383C0C30;
    char_20[9 ]  <=   32'h381C1818;
    char_20[10]  <=   32'h781C1818;
    char_20[11]  <=   32'h781C1808;
    char_20[12]  <=   32'h7C1C300C;
    char_20[13]  <=   32'h381C300C;
    char_20[14]  <=   32'h003C300C;
    char_20[15]  <=   32'h0038300C;
    char_20[16]  <=   32'h0070300C;
    char_20[17]  <=   32'h00F0300C;
    char_20[18]  <=   32'h01E0300C;
    char_20[19]  <=   32'h03C0300C;
    char_20[20]  <=   32'h0780300C;
    char_20[21]  <=   32'h0F00300C;
    char_20[22]  <=   32'h0E061808;
    char_20[23]  <=   32'h1C0E1818;
    char_20[24]  <=   32'h380C1818;
    char_20[25]  <=   32'h701C0C30;
    char_20[26]  <=   32'h7FFC0620;
    char_20[27]  <=   32'h7FFC03C0;
    char_20[28]  <=   32'h00000000;
    char_20[29]  <=   32'h00000000;
    char_20[30]  <=   32'h00000000;
    char_20[31]  <=   32'h00000000;
end 

reg [31:0] char_40[31:0]; 
//40
always @(posedge lcd_pclk) begin
    char_40[0 ]  <=   32'h00000000;
    char_40[1 ]  <=   32'h00000000;
    char_40[2 ]  <=   32'h00000000;
    char_40[3 ]  <=   32'h00000000;
    char_40[4 ]  <=   32'h00000000;
    char_40[5 ]  <=   32'h00000000;
    char_40[6 ]  <=   32'h007003C0;
    char_40[7 ]  <=   32'h00700620;
    char_40[8 ]  <=   32'h00F00C30;
    char_40[9 ]  <=   32'h01F01818;
    char_40[10]  <=   32'h01F01818;
    char_40[11]  <=   32'h03F01808;
    char_40[12]  <=   32'h0370300C;
    char_40[13]  <=   32'h0770300C;
    char_40[14]  <=   32'h0E70300C;
    char_40[15]  <=   32'h0C70300C;
    char_40[16]  <=   32'h1C70300C;
    char_40[17]  <=   32'h1870300C;
    char_40[18]  <=   32'h3870300C;
    char_40[19]  <=   32'h7070300C;
    char_40[20]  <=   32'h6070300C;
    char_40[21]  <=   32'hFFFF300C;
    char_40[22]  <=   32'h00701808;
    char_40[23]  <=   32'h00701818;
    char_40[24]  <=   32'h00701818;
    char_40[25]  <=   32'h00700C30;
    char_40[26]  <=   32'h00F80620;
    char_40[27]  <=   32'h07FE03C0;
    char_40[28]  <=   32'h00000000;
    char_40[29]  <=   32'h00000000;
    char_40[30]  <=   32'h00000000;
    char_40[31]  <=   32'h00000000;
end 
reg [95:0] char_60[31:0]; 
//60/KHZ
always @(posedge lcd_pclk) begin
    char_60[0 ]  <=   96'h000000000000000000000000;
    char_60[1 ]  <=   96'h000000000000000000000000;
    char_60[2 ]  <=   96'h000000000000000000000000;
    char_60[3 ]  <=   96'h000000000002000000000000;
    char_60[4 ]  <=   96'h000000000006000000000000;
    char_60[5 ]  <=   96'h000000000004000000000000;
    char_60[6 ]  <=   96'h03F003C0000C7E7CFC3F1FFE;
    char_60[7 ]  <=   96'h0F38062000081830300C1C0C;
    char_60[8 ]  <=   96'h1E3C0C3000181820300C180C;
    char_60[9 ]  <=   96'h1C3C181800101860300C3018;
    char_60[10]  <=   96'h3818181800301840300C2018;
    char_60[11]  <=   96'h3800180800201880300C0030;
    char_60[12]  <=   96'h7800300C00601880300C0060;
    char_60[13]  <=   96'h7800300C00401900300C0060;
    char_60[14]  <=   96'h7FF0300C00C01900300C00C0;
    char_60[15]  <=   96'h7FF8300C00801B00300C00C0;
    char_60[16]  <=   96'h7C3C300C01801D803FFC0180;
    char_60[17]  <=   96'h781E300C01001D80300C0180;
    char_60[18]  <=   96'h781E300C030018C0300C0300;
    char_60[19]  <=   96'h781E300C020018C0300C0300;
    char_60[20]  <=   96'h781E300C06001860300C0600;
    char_60[21]  <=   96'h781E300C04001860300C0600;
    char_60[22]  <=   96'h781E18080C001830300C0C00;
    char_60[23]  <=   96'h381E181808001830300C1802;
    char_60[24]  <=   96'h3C1C181818001830300C1806;
    char_60[25]  <=   96'h1C1C0C3010001818300C3004;
    char_60[26]  <=   96'h1F78062030001818300C301C;
    char_60[27]  <=   96'h07F003C020007E3EFC3F7FFC;
    char_60[28]  <=   96'h000000006000000000000000;
    char_60[29]  <=   96'h000000004000000000000000;
    char_60[30]  <=   96'h000000000000000000000000;
    char_60[31]  <=   96'h000000000000000000000000;
end 

reg [47:0] char_100[31:0]; 
//100
always @(posedge lcd_pclk) begin
    char_100[0 ]  <=   48'h000000000000;
    char_100[1 ]  <=   48'h000000000000;
    char_100[2 ]  <=   48'h000000000000;
    char_100[3 ]  <=   48'h000000000000;
    char_100[4 ]  <=   48'h000000000000;
    char_100[5 ]  <=   48'h000000000000;
    char_100[6 ]  <=   48'h00C003C003C0;
    char_100[7 ]  <=   48'h03C006200620;
    char_100[8 ]  <=   48'h1FC00C300C30;
    char_100[9 ]  <=   48'h03C018181818;
    char_100[10]  <=   48'h03C018181818;
    char_100[11]  <=   48'h03C018081808;
    char_100[12]  <=   48'h03C0300C300C;
    char_100[13]  <=   48'h03C0300C300C;
    char_100[14]  <=   48'h03C0300C300C;
    char_100[15]  <=   48'h03C0300C300C;
    char_100[16]  <=   48'h03C0300C300C;
    char_100[17]  <=   48'h03C0300C300C;
    char_100[18]  <=   48'h03C0300C300C;
    char_100[19]  <=   48'h03C0300C300C;
    char_100[20]  <=   48'h03C0300C300C;
    char_100[21]  <=   48'h03C0300C300C;
    char_100[22]  <=   48'h03C018081808;
    char_100[23]  <=   48'h03C018181818;
    char_100[24]  <=   48'h03C018181818;
    char_100[25]  <=   48'h03C00C300C30;
    char_100[26]  <=   48'h03E006200620;
    char_100[27]  <=   48'h1FFC03C003C0;
    char_100[28]  <=   48'h000000000000;
    char_100[29]  <=   48'h000000000000;
    char_100[30]  <=   48'h000000000000;
    char_100[31]  <=   48'h000000000000;
end 

reg [47:0] char_150[31:0]; 
//150
always @(posedge lcd_pclk) begin
    char_150[0 ]  <=   48'h000000000000;
    char_150[1 ]  <=   48'h000000000000;
    char_150[2 ]  <=   48'h000000000000;
    char_150[3 ]  <=   48'h000000000000;
    char_150[4 ]  <=   48'h000000000000;
    char_150[5 ]  <=   48'h000000000000;
    char_150[6 ]  <=   48'h00C00FFC03C0;
    char_150[7 ]  <=   48'h03C00FFC0620;
    char_150[8 ]  <=   48'h1FC010000C30;
    char_150[9 ]  <=   48'h03C010001818;
    char_150[10]  <=   48'h03C010001818;
    char_150[11]  <=   48'h03C010001808;
    char_150[12]  <=   48'h03C01000300C;
    char_150[13]  <=   48'h03C01000300C;
    char_150[14]  <=   48'h03C013E0300C;
    char_150[15]  <=   48'h03C01430300C;
    char_150[16]  <=   48'h03C01818300C;
    char_150[17]  <=   48'h03C01008300C;
    char_150[18]  <=   48'h03C0000C300C;
    char_150[19]  <=   48'h03C0000C300C;
    char_150[20]  <=   48'h03C0000C300C;
    char_150[21]  <=   48'h03C0000C300C;
    char_150[22]  <=   48'h03C0300C1808;
    char_150[23]  <=   48'h03C0300C1818;
    char_150[24]  <=   48'h03C020181818;
    char_150[25]  <=   48'h03C020180C30;
    char_150[26]  <=   48'h03E018300620;
    char_150[27]  <=   48'h1FFC07C003C0;
    char_150[28]  <=   48'h000000000000;
    char_150[29]  <=   48'h000000000000;
    char_150[30]  <=   48'h000000000000;
    char_150[31]  <=   48'h000000000000;
end 

reg [47:0] char_200[31:0]; 
//200
always @(posedge lcd_pclk) begin
    char_200[0 ]  <=   48'h000000000000;
    char_200[1 ]  <=   48'h000000000000;
    char_200[2 ]  <=   48'h000000000000;
    char_200[3 ]  <=   48'h000000000000;
    char_200[4 ]  <=   48'h000000000000;
    char_200[5 ]  <=   48'h000000000000;
    char_200[6 ]  <=   48'h0FF003C003C0;
    char_200[7 ]  <=   48'h1E7806200620;
    char_200[8 ]  <=   48'h383C0C300C30;
    char_200[9 ]  <=   48'h381C18181818;
    char_200[10]  <=   48'h781C18181818;
    char_200[11]  <=   48'h781C18081808;
    char_200[12]  <=   48'h7C1C300C300C;
    char_200[13]  <=   48'h381C300C300C;
    char_200[14]  <=   48'h003C300C300C;
    char_200[15]  <=   48'h0038300C300C;
    char_200[16]  <=   48'h0070300C300C;
    char_200[17]  <=   48'h00F0300C300C;
    char_200[18]  <=   48'h01E0300C300C;
    char_200[19]  <=   48'h03C0300C300C;
    char_200[20]  <=   48'h0780300C300C;
    char_200[21]  <=   48'h0F00300C300C;
    char_200[22]  <=   48'h0E0618081808;
    char_200[23]  <=   48'h1C0E18181818;
    char_200[24]  <=   48'h380C18181818;
    char_200[25]  <=   48'h701C0C300C30;
    char_200[26]  <=   48'h7FFC06200620;
    char_200[27]  <=   48'h7FFC03C003C0;
    char_200[28]  <=   48'h000000000000;
    char_200[29]  <=   48'h000000000000;
    char_200[30]  <=   48'h000000000000;
    char_200[31]  <=   48'h000000000000;
end 

reg [63:0] char_x256[31:0]; 
//x256
always @(posedge lcd_pclk) begin
    char_x256[0 ]  <=   64'h0000000000000000;
    char_x256[1 ]  <=   64'h0000000000000000;
    char_x256[2 ]  <=   64'h0000000000000000;
    char_x256[3 ]  <=   64'h0000000000000000;
    char_x256[4 ]  <=   64'h0000000000000000;
    char_x256[5 ]  <=   64'h0000000000000000;
    char_x256[6 ]  <=   64'h000007E00FFC01E0;
    char_x256[7 ]  <=   64'h000008380FFC0618;
    char_x256[8 ]  <=   64'h0000101810000C18;
    char_x256[9 ]  <=   64'h0000200C10000818;
    char_x256[10]  <=   64'h0000200C10001800;
    char_x256[11]  <=   64'h0000300C10001000;
    char_x256[12]  <=   64'h0000300C10001000;
    char_x256[13]  <=   64'h3E7C000C10003000;
    char_x256[14]  <=   64'h0C10001813E033E0;
    char_x256[15]  <=   64'h0E10001814303630;
    char_x256[16]  <=   64'h0620003018183818;
    char_x256[17]  <=   64'h0340006010083808;
    char_x256[18]  <=   64'h034000C0000C300C;
    char_x256[19]  <=   64'h01800180000C300C;
    char_x256[20]  <=   64'h01800300000C300C;
    char_x256[21]  <=   64'h01C00200000C300C;
    char_x256[22]  <=   64'h02600404300C300C;
    char_x256[23]  <=   64'h04600804300C180C;
    char_x256[24]  <=   64'h0430100420181808;
    char_x256[25]  <=   64'h0818200C20180C18;
    char_x256[26]  <=   64'h18183FF818300E30;
    char_x256[27]  <=   64'h7C7E3FF807C003E0;
    char_x256[28]  <=   64'h0000000000000000;
    char_x256[29]  <=   64'h0000000000000000;
    char_x256[30]  <=   64'h0000000000000000;
    char_x256[31]  <=   64'h0000000000000000;
end 
assign   back_en  =  (((pixel_xpos >= PIC_X_START - 1'b1) && (pixel_xpos < PIC_X_START + PIC_WIDTH - 1'b1) && (pixel_ypos >= PIC_Y_START) && (pixel_ypos < PIC_Y_START + PIC_HEIGHT))
                     ||((pixel_xpos >= CHAR_X_START_bx - 1'b1) && (pixel_xpos < CHAR_X_START_bx + CHAR_WIDTH_bx - 1'b1) && (pixel_ypos >= CHAR_Y_START_bx) && (pixel_ypos < CHAR_Y_START_bx + CHAR_HEIGHT))
                     ||((pixel_xpos >= CHAR_X_START_FFT - 1'b1) && (pixel_xpos < CHAR_X_START_FFT + CHAR_WIDTH_FFT - 1'b1) && (pixel_ypos >= CHAR_Y_START_FFT) && (pixel_ypos < CHAR_Y_START_FFT + CHAR_HEIGHT))
                     ||((pixel_xpos >= CHAR_X_START_xsds - 1'b1) && (pixel_xpos < CHAR_X_START_xsds + CHAR_WIDTH_xsds - 1'b1) && (pixel_ypos >= CHAR_Y_START_xsds) && (pixel_ypos < CHAR_Y_START_xsds + CHAR_HEIGHT))
                     ||((pixel_xpos >= CHAR_X_START_ppbj - 1'b1) && (pixel_xpos < CHAR_X_START_ppbj + CHAR_WIDTH_ppbj - 1'b1)&& (pixel_ypos >= CHAR_Y_START_ppbj) && (pixel_ypos < CHAR_Y_START_ppbj + CHAR_HEIGHT)) 
                     ||((pixel_xpos >= CHAR_X_START_sp - 1'b1) && (pixel_xpos < CHAR_X_START_sp + CHAR_WIDTH_sp - 1'b1)&& (pixel_ypos >= CHAR_Y_START_sp) && (pixel_ypos < CHAR_Y_START_sp + CHAR_HEIGHT))
                     ||((pixel_xpos >= CHAR_X_START_fdp - 1'b1) && (pixel_xpos < CHAR_X_START_fdp + CHAR_WIDTH_fdp - 1'b1) && (pixel_ypos >= CHAR_Y_START_fdp) && (pixel_ypos < CHAR_Y_START_fdp + CHAR_HEIGHT)) 
                     ||((pixel_xpos >= CHAR_X_START_0 - 1'b1) && (pixel_xpos < CHAR_X_START_0 + CHAR_WIDTH_0 - 1'b1) && (pixel_ypos >= CHAR_Y_START_0) && (pixel_ypos < CHAR_Y_START_0 + CHAR_HEIGHT))
              //       ||((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1) && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) 
              //       ||((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1) && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT))
              //       ||((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1) && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) 
                     ||((pixel_xpos >= CHAR_X_START_50 - 1'b1) && (pixel_xpos < CHAR_X_START_50 + CHAR_WIDTH_50 - 1'b1) && (pixel_ypos >= CHAR_Y_START_50) && (pixel_ypos < CHAR_Y_START_50 + CHAR_HEIGHT))
                     ||((pixel_xpos >= CHAR_X_START_100 - 1'b1) && (pixel_xpos < CHAR_X_START_100 + CHAR_WIDTH_100 - 1'b1)  && (pixel_ypos >= CHAR_Y_START_100) && (pixel_ypos < CHAR_Y_START_100 + CHAR_HEIGHT))  
                     ||((pixel_xpos >= CHAR_X_START_150 - 1'b1) && (pixel_xpos < CHAR_X_START_150 + CHAR_WIDTH_150 - 1'b1) && (pixel_ypos >= CHAR_Y_START_150) && (pixel_ypos < CHAR_Y_START_150 + CHAR_HEIGHT))
                     ||((pixel_xpos >= CHAR_X_START_200 - 1'b1) && (pixel_xpos < CHAR_X_START_200 + CHAR_WIDTH_200 - 1'b1) && (pixel_ypos >= CHAR_Y_START_200) && (pixel_ypos < CHAR_Y_START_200 + CHAR_HEIGHT))
                     ||((pixel_xpos >= CHAR_X_START_bxzl - 1'b1) && (pixel_xpos < CHAR_X_START_bxzl + CHAR_WIDTH_bxzl - 1'b1) && (pixel_ypos >= CHAR_Y_START_bxzl) && (pixel_ypos < CHAR_Y_START_bxzl + CHAR_HEIGHT))
                     || ((pixel_xpos >= CHAR_X_START_bxpl - 1'b1) && (pixel_xpos < CHAR_X_START_bxpl + CHAR_WIDTH_bxpl - 1'b1) && (pixel_ypos >= CHAR_Y_START_bxpl) && (pixel_ypos < CHAR_Y_START_bxpl + CHAR_HEIGHT))
                     ||((pixel_xpos >= CHAR_X_START_256 - 1'b1) && (pixel_xpos < CHAR_X_START_256 + CHAR_WIDTH_256 - 1'b1) && (pixel_ypos >= CHAR_Y_START_256) && (pixel_ypos < CHAR_Y_START_256 + CHAR_HEIGHT)));



always @(posedge lcd_pclk or negedge rst_n) begin
    if (!rst_n)
        pixel_data <= BACK_COLOR;
    else if( (pixel_xpos >= PIC_X_START - 1'b1) && (pixel_xpos < PIC_X_START + PIC_WIDTH - 1'b1) 
          && (pixel_ypos >= PIC_Y_START) && (pixel_ypos < PIC_Y_START + PIC_HEIGHT) )
        pixel_data <= rom_rd_data ;  //��ʾͼƬ
    else if((pixel_xpos >= CHAR_X_START_bx - 1'b1) && (pixel_xpos < CHAR_X_START_bx + CHAR_WIDTH_bx - 1'b1)
            && (pixel_ypos >= CHAR_Y_START_bx) && (pixel_ypos < CHAR_Y_START_bx + CHAR_HEIGHT)) begin
           if(char_bx[y_cnt_bx][CHAR_WIDTH_bx -1'b1 - x_cnt_bx])
               pixel_data <= CHAR_COLOR;    //��ʾ�ַ� ��ЯƵ����
           else
                   pixel_data <= BLUE;    //��ʾ�ַ�����ı���ɫ
            end   
   else if((pixel_xpos >= CHAR_X_START_bxzl - 1'b1) && (pixel_xpos < CHAR_X_START_bxzl + CHAR_WIDTH_bxzl - 1'b1)
            && (pixel_ypos >= CHAR_Y_START_bxzl) && (pixel_ypos < CHAR_Y_START_bxzl + CHAR_HEIGHT)) begin
           if(char_bxzl[y_cnt_bxzl][CHAR_WIDTH_bxzl -1'b1 - x_cnt_bxzl])
               pixel_data <= CHAR_COLOR;    //��ʾ�ַ� �������ࣺ
           else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
            end   
    else if((pixel_xpos >= CHAR_X_START_bxpl - 1'b1) && (pixel_xpos < CHAR_X_START_bxpl + CHAR_WIDTH_bxpl - 1'b1)
                && (pixel_ypos >= CHAR_Y_START_bxpl) && (pixel_ypos < CHAR_Y_START_bxpl + CHAR_HEIGHT)) begin
               if(char_bxpl[y_cnt_bxpl][CHAR_WIDTH_bxpl -1'b1 - x_cnt_bxpl])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� ����Ƶ�ʣ�
               else
                       pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
                end           
    else if((pixel_xpos >= CHAR_X_START_FFT - 1'b1) && (pixel_xpos < CHAR_X_START_FFT + CHAR_WIDTH_FFT - 1'b1)
                && (pixel_ypos >= CHAR_Y_START_FFT) && (pixel_ypos < CHAR_Y_START_FFT + CHAR_HEIGHT)) begin
         if(char_FFT[y_cnt_FFT][CHAR_WIDTH_FFT -1'b1 - x_cnt_FFT])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� FFT:256
         else
                       pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
                end
   else if((pixel_xpos >= CHAR_X_START_xsds - 1'b1) && (pixel_xpos < CHAR_X_START_xsds + CHAR_WIDTH_xsds - 1'b1)
                    && (pixel_ypos >= CHAR_Y_START_xsds) && (pixel_ypos < CHAR_Y_START_xsds + CHAR_HEIGHT)) begin
        if(char_xsds[y_cnt_xsds][CHAR_WIDTH_xsds -1'b1 - x_cnt_xsds])
                pixel_data <= CHAR_COLOR;    //��ʾ�ַ� ��ʾ������128
        else
                pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_ppbj - 1'b1) && (pixel_xpos < CHAR_X_START_ppbj + CHAR_WIDTH_ppbj - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_ppbj) && (pixel_ypos < CHAR_Y_START_ppbj + CHAR_HEIGHT)) begin
            if(char_ppbj[y_cnt_ppbj][CHAR_WIDTH_ppbj -1'b1 - x_cnt_ppbj])
                    pixel_data <= CHAR_COLOR;    //��ʾ�ַ� Ƶ�ײ�����5
     else
                    pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
      end
      else if((pixel_xpos >= CHAR_X_START_sp - 1'b1) && (pixel_xpos < CHAR_X_START_sp + CHAR_WIDTH_sp - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_sp) && (pixel_ypos < CHAR_Y_START_sp + CHAR_HEIGHT)) begin
                if(char_sp[y_cnt_sp][CHAR_WIDTH_sp -1'b1 - x_cnt_sp])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� ˮƽ��20/div
     else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_fdp - 1'b1) && (pixel_xpos < CHAR_X_START_fdp + CHAR_WIDTH_fdp - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_fdp) && (pixel_ypos < CHAR_Y_START_fdp + CHAR_HEIGHT)) begin
                if(char_fdp[y_cnt_fdp][CHAR_WIDTH_fdp -1'b1 - x_cnt_fdp])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� ������
     else
                   pixel_data <= BLUE;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_0 - 1'b1) && (pixel_xpos < CHAR_X_START_0 + CHAR_WIDTH_0 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_0) && (pixel_ypos < CHAR_Y_START_0 + CHAR_HEIGHT)) begin
                if(char_0[y_cnt_0][CHAR_WIDTH_0 -1'b1 - x_cnt_0])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� 0
     else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
                if(char_20[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� 20
     else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                if(char_40[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� 40
     else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                if(char_60[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� 60/KHZ
     else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_50 - 1'b1) && (pixel_xpos < CHAR_X_START_50 + CHAR_WIDTH_50 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_50) && (pixel_ypos < CHAR_Y_START_50 + CHAR_HEIGHT)) begin
                if(char_50[y_cnt_50][CHAR_WIDTH_50 -1'b1 - x_cnt_50])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� 50
     else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_100 - 1'b1) && (pixel_xpos < CHAR_X_START_100 + CHAR_WIDTH_100 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_100) && (pixel_ypos < CHAR_Y_START_100 + CHAR_HEIGHT)) begin
                if(char_100[y_cnt_100][CHAR_WIDTH_100 -1'b1 - x_cnt_100])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� 100
     else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_150 - 1'b1) && (pixel_xpos < CHAR_X_START_150 + CHAR_WIDTH_150 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_150) && (pixel_ypos < CHAR_Y_START_150 + CHAR_HEIGHT)) begin
                if(char_150[y_cnt_150][CHAR_WIDTH_150 -1'b1 - x_cnt_150])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� 150
     else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_200 - 1'b1) && (pixel_xpos < CHAR_X_START_200 + CHAR_WIDTH_200 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_200) && (pixel_ypos < CHAR_Y_START_200 + CHAR_HEIGHT)) begin
                if(char_200[y_cnt_200][CHAR_WIDTH_200 -1'b1 - x_cnt_200])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� 200
     else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
     else if((pixel_xpos >= CHAR_X_START_256 - 1'b1) && (pixel_xpos < CHAR_X_START_256 + CHAR_WIDTH_256 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_256) && (pixel_ypos < CHAR_Y_START_256 + CHAR_HEIGHT)) begin
                if(char_x256[y_cnt_256][CHAR_WIDTH_256 -1'b1 - x_cnt_256])
                   pixel_data <= CHAR_COLOR;    //��ʾ�ַ� x256
     else
                   pixel_data <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
     end
    else 
        pixel_data <= BACK_COLOR;
    end 
//���ݵ�ǰɨ���ĺ�������ΪROM��ַ��ֵ
always @(posedge lcd_pclk or negedge rst_n) begin
    if(!rst_n)
        rom_addr <= 11'd0;
    //����������λ��ͼƬ��ʾ����ʱ,�ۼ�ROM��ַ    
    else if((pixel_ypos >= PIC_Y_START) && (pixel_ypos < PIC_Y_START + PIC_HEIGHT) 
        && (pixel_xpos >= PIC_X_START - 2'd2) && (pixel_xpos < PIC_X_START + PIC_WIDTH - 2'd2)) 
        rom_addr <= rom_addr + 1'b1;
    //����������λ��ͼƬ�������һ�����ص�ʱ,ROM��ַ����    
    else if((pixel_ypos >= PIC_Y_START + PIC_HEIGHT))
        rom_addr <= 11'd0;
end

assign wave_en = ((pixel_xpos >= CHAR_X_START_zxb - 1'b1) && (pixel_xpos < CHAR_X_START_zxb + CHAR_WIDTH_zxb - 1'b1)&& (pixel_ypos >= CHAR_Y_START_zxb) && (pixel_ypos < CHAR_Y_START_zxb + CHAR_HEIGHT));
always @(posedge lcd_pclk or negedge rst_n) begin
    if (!rst_n)
        pixel_data_wave <= BACK_COLOR;
    else case(wave_choose)
    2'b00: if((pixel_xpos >= CHAR_X_START_zxb - 1'b1) && (pixel_xpos < CHAR_X_START_zxb + CHAR_WIDTH_zxb - 1'b1)
            && (pixel_ypos >= CHAR_Y_START_zxb) && (pixel_ypos < CHAR_Y_START_zxb + CHAR_HEIGHT)) begin
           if(char_zxb[y_cnt_zxb][CHAR_WIDTH_zxb -1'b1 - x_cnt_zxb])
               pixel_data_wave <= CHAR_COLOR;    //��ʾ�ַ� 
           else
                   pixel_data_wave <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
            end   
            else
                pixel_data_wave <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
    2'b01:if((pixel_xpos >= CHAR_X_START_sjb - 1'b1) && (pixel_xpos < CHAR_X_START_sjb + CHAR_WIDTH_sjb - 1'b1)
                && (pixel_ypos >= CHAR_Y_START_sjb) && (pixel_ypos < CHAR_Y_START_sjb + CHAR_HEIGHT)) begin
         if(char_sjb[y_cnt_sjb][CHAR_WIDTH_sjb -1'b1 - x_cnt_sjb])
                   pixel_data_wave <= CHAR_COLOR;    //��ʾ�ַ� 
         else
                       pixel_data_wave <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
                end
         else
                    pixel_data_wave <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
    2'b10: if((pixel_xpos >= CHAR_X_START_jcb - 1'b1) && (pixel_xpos < CHAR_X_START_jcb + CHAR_WIDTH_jcb - 1'b1)
                    && (pixel_ypos >= CHAR_Y_START_jcb) && (pixel_ypos < CHAR_Y_START_jcb + CHAR_HEIGHT)) begin
                   if(char_jcb[y_cnt_jcb][CHAR_WIDTH_jcb -1'b1 - x_cnt_jcb])
                       pixel_data_wave <= CHAR_COLOR;    //��ʾ�ַ� 
                   else
                           pixel_data_wave <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
                    end   
                    else
                        pixel_data_wave <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
    2'b11:if((pixel_xpos >= CHAR_X_START_fb - 1'b1) && (pixel_xpos < CHAR_X_START_fb + CHAR_WIDTH_fb - 1'b1)
                        && (pixel_ypos >= CHAR_Y_START_fb) && (pixel_ypos < CHAR_Y_START_fb + CHAR_HEIGHT)) begin
                 if(char_fb[y_cnt_fb][CHAR_WIDTH_fb -1'b1 - x_cnt_fb])
                           pixel_data_wave <= CHAR_COLOR;    //��ʾ�ַ� 
                 else
                               pixel_data_wave <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
                        end
                 else
                            pixel_data_wave <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
    default: if((pixel_xpos >= CHAR_X_START_fb - 1'b1) && (pixel_xpos < CHAR_X_START_fb + CHAR_WIDTH_fb - 1'b1)
                 && (pixel_ypos >= CHAR_Y_START_fb) && (pixel_ypos < CHAR_Y_START_fb + CHAR_HEIGHT)) begin
           if(char_fb[y_cnt_fb][CHAR_WIDTH_fb -1'b1 - x_cnt_fb])
                               pixel_data_wave <= CHAR_COLOR;    //��ʾ�ַ� 
                else
                               pixel_data_wave <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
                   end
                  else
                            pixel_data_wave <= BACK_COLOR;    //��ʾ�ַ�����ı���ɫ
    endcase
end 
//ROM���洢ͼƬ
ziguanrom1 ziguanrom1_isnt (
  .addr(rom_addr),          // input [10:0]
  .clk(lcd_pclk),            // input
  .rst(~rst_n),            // input
  .rd_data(rom_rd_data)     // output [23:0]
);

endmodule 







