module fft_div_adaptive(
    input             lcd_pclk  ,               //lcd驱动时钟
    input             sys_rst_n ,               //复位信号
	input      [35:0] data_d0      ,
    input      [10:0] pixel_xpos,               //像素点横坐标   在例化时将低位宽的像素坐标拼接0即可满足该模块的位宽
    input      [10:0] pixel_ypos,               //像素点纵坐标
    input      [11:0] freq_adj,
    output            fre_eq_diven,
    output reg [23:0] pixel_data                //像素点数据

   );

   localparam BACK_COLOR  = 24'hffffff; //背景色，白色
   //localparam CHAR_COLOR  = 24'hff0000; //字符颜色，红色
   localparam BLUE   = 24'b00000000_00000000_11111111;     //RGB888 蓝色
   localparam CHAR_COLOR  = 24'b00000000_00000000_00000000; //字符颜色，黑色


   localparam CHAR_HEIGHT = 11'd32;     //字符高度
   localparam CHAR_X_START_680= 11'd224;     //字符起始点横坐标 20   32x32
   localparam CHAR_Y_START_680= 11'd438;    //字符起始点纵坐标    保持三位宽  少于的补上空格
   localparam CHAR_WIDTH_680 = 11'd64;    //字符宽度, 
   wire  [10:0]  x_cnt_680;       //横坐标计数器
   wire  [10:0]  y_cnt_680;       //纵坐标计数器
   assign  x_cnt_680 = pixel_xpos + 1'b1  - CHAR_X_START_680; //像素点相对于字符区域起始点水平坐标
   assign  y_cnt_680 = pixel_ypos - CHAR_Y_START_680; //像素点相对于字符区域起始点垂直坐标
   
   localparam CHAR_X_START_135= 11'd424;     //字符起始点横坐标 40   32x32
   localparam CHAR_Y_START_135= 11'd438;    //字符起始点纵坐标 
   localparam CHAR_WIDTH_135 = 11'd64;    //字符宽度, 
   wire  [10:0]  x_cnt_135;       //横坐标计数器
   wire  [10:0]  y_cnt_135;       //纵坐标计数器
   assign  x_cnt_135 = pixel_xpos + 1'b1  - CHAR_X_START_135; //像素点相对于字符区域起始点水平坐标
   assign  y_cnt_135 = pixel_ypos - CHAR_Y_START_135; //像素点相对于字符区域起始点垂直坐标
   


   localparam CHAR_X_START_20= 11'd232;     //字符起始点横坐标 20   32x32
   localparam CHAR_Y_START_20= 11'd438;    //字符起始点纵坐标    保持三位宽  少于的补上空格
   localparam CHAR_WIDTH_20  = 11'd48;    //字符宽度, 
   wire  [10:0]  x_cnt_20;       //横坐标计数器
   wire  [10:0]  y_cnt_20;       //纵坐标计数器
   assign  x_cnt_20 = pixel_xpos + 1'b1  - CHAR_X_START_20; //像素点相对于字符区域起始点水平坐标
   assign  y_cnt_20 = pixel_ypos - CHAR_Y_START_20; //像素点相对于字符区域起始点垂直坐标
   
   localparam CHAR_X_START_40= 11'd432;     //字符起始点横坐标 40   32x32
   localparam CHAR_Y_START_40= 11'd438;    //字符起始点纵坐标 
   localparam CHAR_WIDTH_40  = 11'd48;    //字符宽度, 
   wire  [10:0]  x_cnt_40;       //横坐标计数器
   wire  [10:0]  y_cnt_40;       //纵坐标计数器
   assign  x_cnt_40 = pixel_xpos + 1'b1  - CHAR_X_START_40; //像素点相对于字符区域起始点水平坐标
   assign  y_cnt_40 = pixel_ypos - CHAR_Y_START_40; //像素点相对于字符区域起始点垂直坐标
   
   localparam CHAR_X_START_60= 11'd632;     //字符起始点横坐标 60/KHZ   96x32
   localparam CHAR_Y_START_60= 11'd438;    //字符起始点纵坐标 
   localparam CHAR_WIDTH_60  = 11'd112;    //字符宽度, 
   wire  [10:0]  x_cnt_60;       //横坐标计数器
   wire  [10:0]  y_cnt_60;       //纵坐标计数器
   assign  x_cnt_60 = pixel_xpos + 1'b1  - CHAR_X_START_60; //像素点相对于字符区域起始点水平坐标
   assign  y_cnt_60 = pixel_ypos - CHAR_Y_START_60; //像素点相对于字符区域起始点垂直坐标


   localparam CHAR_X_START_1000= 11'd616;     //字符起始点横坐标 60/KHZ   96x32
   localparam CHAR_Y_START_1000= 11'd438;    //字符起始点纵坐标 
   localparam CHAR_WIDTH_1000 = 11'd128;    //字符宽度, 
   wire  [10:0]  x_cnt_1000;       //横坐标计数器
   wire  [10:0]  y_cnt_1000;       //纵坐标计数器
   assign  x_cnt_1000 = pixel_xpos + 1'b1  - CHAR_X_START_1000; //像素点相对于字符区域起始点水平坐标
   assign  y_cnt_1000 = pixel_ypos - CHAR_Y_START_1000; //像素点相对于字符区域起始点垂直坐标
   
assign  fre_eq_diven  = (((pixel_xpos >= CHAR_X_START_1000 - 1'b1) && (pixel_xpos < CHAR_X_START_1000 + CHAR_WIDTH_1000 - 1'b1) && (pixel_ypos >= CHAR_Y_START_1000) && (pixel_ypos < CHAR_Y_START_1000 + CHAR_HEIGHT))
                        ||((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1) && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) 
                        ||((pixel_xpos >= CHAR_X_START_680 - 1'b1) && (pixel_xpos < CHAR_X_START_680 + CHAR_WIDTH_680 - 1'b1) && (pixel_ypos >= CHAR_Y_START_680) && (pixel_ypos < CHAR_Y_START_680 + CHAR_HEIGHT)) 
                        ||((pixel_xpos >= CHAR_X_START_135 - 1'b1) && (pixel_xpos < CHAR_X_START_135 + CHAR_WIDTH_135 - 1'b1) && (pixel_ypos >= CHAR_Y_START_135) && (pixel_ypos < CHAR_Y_START_135 + CHAR_HEIGHT))
                        ||((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1) && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT))
                        ||((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1) && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) );


 reg [47:0] char_1d3 [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_1d3[0 ]  <=   48'h000000000000;
                            char_1d3[1 ]  <=   48'h000000000000;
                            char_1d3[2 ]  <=   48'h000000000000;
                            char_1d3[3 ]  <=   48'h000000000000;
                            char_1d3[4 ]  <=   48'h000000000000;
                            char_1d3[5 ]  <=   48'h000000000000;
                            char_1d3[6 ]  <=   48'h00C0000007C0;
                            char_1d3[7 ]  <=   48'h03C000001860;
                            char_1d3[8 ]  <=   48'h1FC000003030;
                            char_1d3[9 ]  <=   48'h03C000003018;
                            char_1d3[10]  <=   48'h03C000003018;
                            char_1d3[11]  <=   48'h03C000003018;
                            char_1d3[12]  <=   48'h03C000000018;
                            char_1d3[13]  <=   48'h03C000000018;
                            char_1d3[14]  <=   48'h03C000000030;
                            char_1d3[15]  <=   48'h03C000000060;
                            char_1d3[16]  <=   48'h03C0000003C0;
                            char_1d3[17]  <=   48'h03C000000070;
                            char_1d3[18]  <=   48'h03C000000018;
                            char_1d3[19]  <=   48'h03C000000008;
                            char_1d3[20]  <=   48'h03C00000000C;
                            char_1d3[21]  <=   48'h03C00000000C;
                            char_1d3[22]  <=   48'h03C00000300C;
                            char_1d3[23]  <=   48'h03C00000300C;
                            char_1d3[24]  <=   48'h03C018003008;
                            char_1d3[25]  <=   48'h03C03C003018;
                            char_1d3[26]  <=   48'h03E03C001830;
                            char_1d3[27]  <=   48'h1FFC180007C0;
                            char_1d3[28]  <=   48'h000000000000;
                            char_1d3[29]  <=   48'h000000000000;
                            char_1d3[30]  <=   48'h000000000000;
                            char_1d3[31]  <=   48'h000000000000;
end 

reg [47:0] char_640 [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_640[0 ]  <=   48'h000000000000;
                            char_640[1 ]  <=   48'h000000000000;
                            char_640[2 ]  <=   48'h000000000000;
                            char_640[3 ]  <=   48'h000000000000;
                            char_640[4 ]  <=   48'h000000000000;
                            char_640[5 ]  <=   48'h000000000000;
                            char_640[6 ]  <=   48'h03F0006003C0;
                            char_640[7 ]  <=   48'h0F3800600620;
                            char_640[8 ]  <=   48'h1E3C00E00C30;
                            char_640[9 ]  <=   48'h1C3C00E01818;
                            char_640[10]  <=   48'h381801601818;
                            char_640[11]  <=   48'h380001601808;
                            char_640[12]  <=   48'h78000260300C;
                            char_640[13]  <=   48'h78000460300C;
                            char_640[14]  <=   48'h7FF00460300C;
                            char_640[15]  <=   48'h7FF80860300C;
                            char_640[16]  <=   48'h7C3C0860300C;
                            char_640[17]  <=   48'h781E1060300C;
                            char_640[18]  <=   48'h781E3060300C;
                            char_640[19]  <=   48'h781E2060300C;
                            char_640[20]  <=   48'h781E4060300C;
                            char_640[21]  <=   48'h781E7FFC300C;
                            char_640[22]  <=   48'h781E00601808;
                            char_640[23]  <=   48'h381E00601818;
                            char_640[24]  <=   48'h3C1C00601818;
                            char_640[25]  <=   48'h1C1C00600C30;
                            char_640[26]  <=   48'h1F7800600620;
                            char_640[27]  <=   48'h07F003FC03C0;
                            char_640[28]  <=   48'h000000000000;
                            char_640[29]  <=   48'h000000000000;
                            char_640[30]  <=   48'h000000000000;
                            char_640[31]  <=   48'h000000000000;
end 



                        reg [47:0] char_2d5 [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_2d5[0 ]  <=   48'h000000000000;
                            char_2d5[1 ]  <=   48'h000000000000;
                            char_2d5[2 ]  <=   48'h000000000000;
                            char_2d5[3 ]  <=   48'h000000000000;
                            char_2d5[4 ]  <=   48'h000000000000;
                            char_2d5[5 ]  <=   48'h000000000000;
                            char_2d5[6 ]  <=   48'h07E000000FFC;
                            char_2d5[7 ]  <=   48'h083800000FFC;
                            char_2d5[8 ]  <=   48'h101800001000;
                            char_2d5[9 ]  <=   48'h200C00001000;
                            char_2d5[10]  <=   48'h200C00001000;
                            char_2d5[11]  <=   48'h300C00001000;
                            char_2d5[12]  <=   48'h300C00001000;
                            char_2d5[13]  <=   48'h000C00001000;
                            char_2d5[14]  <=   48'h0018000013E0;
                            char_2d5[15]  <=   48'h001800001430;
                            char_2d5[16]  <=   48'h003000001818;
                            char_2d5[17]  <=   48'h006000001008;
                            char_2d5[18]  <=   48'h00C00000000C;
                            char_2d5[19]  <=   48'h01800000000C;
                            char_2d5[20]  <=   48'h03000000000C;
                            char_2d5[21]  <=   48'h02000000000C;
                            char_2d5[22]  <=   48'h04040000300C;
                            char_2d5[23]  <=   48'h08040000300C;
                            char_2d5[24]  <=   48'h100418002018;
                            char_2d5[25]  <=   48'h200C3C002018;
                            char_2d5[26]  <=   48'h3FF83C001830;
                            char_2d5[27]  <=   48'h3FF8180007C0;
                            char_2d5[28]  <=   48'h000000000000;
                            char_2d5[29]  <=   48'h000000000000;
                            char_2d5[30]  <=   48'h000000000000;
                            char_2d5[31]  <=   48'h000000000000;
end 

reg [111:0] char_3d8mhz [31:0];
//空2空 对应MHZ级别
   always @(posedge lcd_pclk) begin
    char_3d8mhz[0 ]  <=   112'h0000000000000000000000000000;
    char_3d8mhz[1 ]  <=   112'h0000000000000000000000000000;
    char_3d8mhz[2 ]  <=   112'h0000000000000000000000000000;
    char_3d8mhz[3 ]  <=   112'h0000000000000002000000000000;
    char_3d8mhz[4 ]  <=   112'h0000000000000006000000000000;
    char_3d8mhz[5 ]  <=   112'h0000000000000004000000000000;
    char_3d8mhz[6 ]  <=   112'h0FE0000007E0000CF00FFC3F1FFE;
    char_3d8mhz[7 ]  <=   112'h1CF000000C300008381C300C1C0C;
    char_3d8mhz[8 ]  <=   112'h3878000018180018381C300C180C;
    char_3d8mhz[9 ]  <=   112'h383C0000300C0010381C300C3018;
    char_3d8mhz[10]  <=   112'h383C0000300C0030381C300C2018;
    char_3d8mhz[11]  <=   112'h383C0000300C0020382C300C0030;
    char_3d8mhz[12]  <=   112'h003C0000380C00602C2C300C0060;
    char_3d8mhz[13]  <=   112'h00380000380800402C2C300C0060;
    char_3d8mhz[14]  <=   112'h007800001E1800C02C2C300C00C0;
    char_3d8mhz[15]  <=   112'h01F000000F2000802C4C300C00C0;
    char_3d8mhz[16]  <=   112'h07E0000007C001802C4C3FFC0180;
    char_3d8mhz[17]  <=   112'h00F8000018F00100264C300C0180;
    char_3d8mhz[18]  <=   112'h0038000030780300264C300C0300;
    char_3d8mhz[19]  <=   112'h001C000030380200264C300C0300;
    char_3d8mhz[20]  <=   112'h001E0000601C0600268C300C0600;
    char_3d8mhz[21]  <=   112'h001E0000600C0400228C300C0600;
    char_3d8mhz[22]  <=   112'h381E0000600C0C00238C300C0C00;
    char_3d8mhz[23]  <=   112'h781E0000600C0800238C300C1802;
    char_3d8mhz[24]  <=   112'h781C1800600C1800230C300C1806;
    char_3d8mhz[25]  <=   112'h383C3C0030181000230C300C3004;
    char_3d8mhz[26]  <=   112'h3CF83C0018303000210C300C301C;
    char_3d8mhz[27]  <=   112'h0FE0180007C02000F13FFC3F7FFC;
    char_3d8mhz[28]  <=   112'h0000000000006000000000000000;
    char_3d8mhz[29]  <=   112'h0000000000004000000000000000;
    char_3d8mhz[30]  <=   112'h0000000000000000000000000000;
    char_3d8mhz[31]  <=   112'h0000000000000000000000000000;
end 

reg [111:0] char_7d6mhz [31:0];
//空2空 对应MHZ级别
   always @(posedge lcd_pclk) begin
    char_7d6mhz[0 ]  <=   112'h0000000000000000000000000000;
    char_7d6mhz[1 ]  <=   112'h0000000000000000000000000000;
    char_7d6mhz[2 ]  <=   112'h0000000000000000000000000000;
    char_7d6mhz[3 ]  <=   112'h0000000000000002000000000000;
    char_7d6mhz[4 ]  <=   112'h0000000000000006000000000000;
    char_7d6mhz[5 ]  <=   112'h0000000000000004000000000000;
    char_7d6mhz[6 ]  <=   112'h3FFE000001E0000CF00FFC3F1FFE;
    char_7d6mhz[7 ]  <=   112'h3FFE000006180008381C300C1C0C;
    char_7d6mhz[8 ]  <=   112'h381C00000C180018381C300C180C;
    char_7d6mhz[9 ]  <=   112'h3018000008180010381C300C3018;
    char_7d6mhz[10]  <=   112'h7038000018000030381C300C2018;
    char_7d6mhz[11]  <=   112'h2030000010000020382C300C0030;
    char_7d6mhz[12]  <=   112'h00700000100000602C2C300C0060;
    char_7d6mhz[13]  <=   112'h00600000300000402C2C300C0060;
    char_7d6mhz[14]  <=   112'h00E0000033E000C02C2C300C00C0;
    char_7d6mhz[15]  <=   112'h00E00000363000802C4C300C00C0;
    char_7d6mhz[16]  <=   112'h01C00000381801802C4C3FFC0180;
    char_7d6mhz[17]  <=   112'h01C0000038080100264C300C0180;
    char_7d6mhz[18]  <=   112'h03C00000300C0300264C300C0300;
    char_7d6mhz[19]  <=   112'h03800000300C0200264C300C0300;
    char_7d6mhz[20]  <=   112'h03800000300C0600268C300C0600;
    char_7d6mhz[21]  <=   112'h03800000300C0400228C300C0600;
    char_7d6mhz[22]  <=   112'h07800000300C0C00238C300C0C00;
    char_7d6mhz[23]  <=   112'h07800000180C0800238C300C1802;
    char_7d6mhz[24]  <=   112'h0780180018081800230C300C1806;
    char_7d6mhz[25]  <=   112'h07803C000C181000230C300C3004;
    char_7d6mhz[26]  <=   112'h07803C000E303000210C300C301C;
    char_7d6mhz[27]  <=   112'h0780180003E02000F13FFC3F7FFC;
    char_7d6mhz[28]  <=   112'h0000000000006000000000000000;
    char_7d6mhz[29]  <=   112'h0000000000004000000000000000;
    char_7d6mhz[30]  <=   112'h0000000000000000000000000000;
    char_7d6mhz[31]  <=   112'h0000000000000000000000000000;
end 
                            
reg [111:0] char_15mhz [31:0];
//空2空 对应MHZ级别
   always @(posedge lcd_pclk) begin
    char_15mhz[0 ]  <=   112'h0000000000000000000000000000;
    char_15mhz[1 ]  <=   112'h0000000000000000000000000000;
    char_15mhz[2 ]  <=   112'h0000000000000000000000000000;
    char_15mhz[3 ]  <=   112'h0000000000000002000000000000;
    char_15mhz[4 ]  <=   112'h0000000000000006000000000000;
    char_15mhz[5 ]  <=   112'h0000000000000004000000000000;
    char_15mhz[6 ]  <=   112'h000000800FFC000CF00FFC3F1FFE;
    char_15mhz[7 ]  <=   112'h000001800FFC0008381C300C1C0C;
    char_15mhz[8 ]  <=   112'h00001F8010000018381C300C180C;
    char_15mhz[9 ]  <=   112'h0000018010000010381C300C3018;
    char_15mhz[10]  <=   112'h0000018010000030381C300C2018;
    char_15mhz[11]  <=   112'h0000018010000020382C300C0030;
    char_15mhz[12]  <=   112'h00000180100000602C2C300C0060;
    char_15mhz[13]  <=   112'h00000180100000402C2C300C0060;
    char_15mhz[14]  <=   112'h0000018013E000C02C2C300C00C0;
    char_15mhz[15]  <=   112'h00000180143000802C4C300C00C0;
    char_15mhz[16]  <=   112'h00000180181801802C4C3FFC0180;
    char_15mhz[17]  <=   112'h0000018010080100264C300C0180;
    char_15mhz[18]  <=   112'h00000180000C0300264C300C0300;
    char_15mhz[19]  <=   112'h00000180000C0200264C300C0300;
    char_15mhz[20]  <=   112'h00000180000C0600268C300C0600;
    char_15mhz[21]  <=   112'h00000180000C0400228C300C0600;
    char_15mhz[22]  <=   112'h00000180300C0C00238C300C0C00;
    char_15mhz[23]  <=   112'h00000180300C0800238C300C1802;
    char_15mhz[24]  <=   112'h0000018020181800230C300C1806;
    char_15mhz[25]  <=   112'h0000018020181000230C300C3004;
    char_15mhz[26]  <=   112'h000003C018303000210C300C301C;
    char_15mhz[27]  <=   112'h00001FF807C02000F13FFC3F7FFC;
    char_15mhz[28]  <=   112'h0000000000006000000000000000;
    char_15mhz[29]  <=   112'h0000000000004000000000000000;
    char_15mhz[30]  <=   112'h0000000000000000000000000000;
    char_15mhz[31]  <=   112'h0000000000000000000000000000;  
end 
                    
reg [111:0] char_960khz [31:0];
//空2空 对应MHZ级别
   always @(posedge lcd_pclk) begin
    char_960khz[0 ]  <=   112'h0000000000000000000000000000;
    char_960khz[1 ]  <=   112'h0000000000000000000000000000;
    char_960khz[2 ]  <=   112'h0000000000000000000000000000;
    char_960khz[3 ]  <=   112'h0000000000000002000000000000;
    char_960khz[4 ]  <=   112'h0000000000000006000000000000;
    char_960khz[5 ]  <=   112'h0000000000000004000000000000;
    char_960khz[6 ]  <=   112'h0FE001E003C0000C7E7CFC3F1FFE;
    char_960khz[7 ]  <=   112'h1EF00618062000081830300C1C0C;
    char_960khz[8 ]  <=   112'h38380C180C3000181820300C180C;
    char_960khz[9 ]  <=   112'h783C0818181800101860300C3018;
    char_960khz[10]  <=   112'h781C1800181800301840300C2018;
    char_960khz[11]  <=   112'h701E1000180800201880300C0030;
    char_960khz[12]  <=   112'h701E1000300C00601880300C0060;
    char_960khz[13]  <=   112'h701E3000300C00401900300C0060;
    char_960khz[14]  <=   112'h701E33E0300C00C01900300C00C0;
    char_960khz[15]  <=   112'h781E3630300C00801B00300C00C0;
    char_960khz[16]  <=   112'h783E3818300C01801D803FFC0180;
    char_960khz[17]  <=   112'h787E3808300C01001D80300C0180;
    char_960khz[18]  <=   112'h3FFE300C300C030018C0300C0300;
    char_960khz[19]  <=   112'h1FDE300C300C020018C0300C0300;
    char_960khz[20]  <=   112'h001E300C300C06001860300C0600;
    char_960khz[21]  <=   112'h001C300C300C04001860300C0600;
    char_960khz[22]  <=   112'h003C300C18080C001830300C0C00;
    char_960khz[23]  <=   112'h1838180C181808001830300C1802;
    char_960khz[24]  <=   112'h3C381808181818001830300C1806;
    char_960khz[25]  <=   112'h3C700C180C3010001818300C3004;
    char_960khz[26]  <=   112'h3DE00E30062030001818300C301C;
    char_960khz[27]  <=   112'h1FC003E003C020007E3EFC3F7FFC;
    char_960khz[28]  <=   112'h0000000000006000000000000000;
    char_960khz[29]  <=   112'h0000000000004000000000000000;
    char_960khz[30]  <=   112'h0000000000000000000000000000;
    char_960khz[31]  <=   112'h0000000000000000000000000000;  
end 
              
reg [63:0] char_1270 [31:0];
//空2空 对应MHZ级别
   always @(posedge lcd_pclk) begin
    char_1270[0 ]  <=   64'h0000000000000000;
    char_1270[1 ]  <=   64'h0000000000000000;
    char_1270[2 ]  <=   64'h0000000000000000;
    char_1270[3 ]  <=   64'h0000000000000000;
    char_1270[4 ]  <=   64'h0000000000000000;
    char_1270[5 ]  <=   64'h0000000000000000;
    char_1270[6 ]  <=   64'h00C007E01FFC03C0;
    char_1270[7 ]  <=   64'h03C008381FFC0620;
    char_1270[8 ]  <=   64'h1FC0101810080C30;
    char_1270[9 ]  <=   64'h03C0200C30101818;
    char_1270[10]  <=   64'h03C0200C20101818;
    char_1270[11]  <=   64'h03C0300C20201808;
    char_1270[12]  <=   64'h03C0300C0020300C;
    char_1270[13]  <=   64'h03C0000C0040300C;
    char_1270[14]  <=   64'h03C000180040300C;
    char_1270[15]  <=   64'h03C000180040300C;
    char_1270[16]  <=   64'h03C000300080300C;
    char_1270[17]  <=   64'h03C000600080300C;
    char_1270[18]  <=   64'h03C000C00100300C;
    char_1270[19]  <=   64'h03C001800100300C;
    char_1270[20]  <=   64'h03C003000100300C;
    char_1270[21]  <=   64'h03C002000100300C;
    char_1270[22]  <=   64'h03C0040403001808;
    char_1270[23]  <=   64'h03C0080403001818;
    char_1270[24]  <=   64'h03C0100403001818;
    char_1270[25]  <=   64'h03C0200C03000C30;
    char_1270[26]  <=   64'h03E03FF803000620;
    char_1270[27]  <=   64'h1FFC3FF8030003C0;
    char_1270[28]  <=   64'h0000000000000000;
    char_1270[29]  <=   64'h0000000000000000;
    char_1270[30]  <=   64'h0000000000000000;
    char_1270[31]  <=   64'h0000000000000000; 
end 


reg [127:0] char_1900khz [31:0];
//空2空 对应MHZ级别
   always @(posedge lcd_pclk) begin
    char_1900khz[0 ]  <=   128'h00000000000000000000000000000000;
    char_1900khz[1 ]  <=   128'h00000000000000000000000000000000;
    char_1900khz[2 ]  <=   128'h00000000000000000000000000000000;
    char_1900khz[3 ]  <=   128'h00000000000000000002000000000000;
    char_1900khz[4 ]  <=   128'h00000000000000000006000000000000;
    char_1900khz[5 ]  <=   128'h00000000000000000004000000000000;
    char_1900khz[6 ]  <=   128'h00C007C003C003C0000C7E7CFC3F1FFE;
    char_1900khz[7 ]  <=   128'h03C018200620062000081830300C1C0C;
    char_1900khz[8 ]  <=   128'h1FC030100C300C3000181820300C180C;
    char_1900khz[9 ]  <=   128'h03C030181818181800101860300C3018;
    char_1900khz[10]  <=   128'h03C060081818181800301840300C2018;
    char_1900khz[11]  <=   128'h03C0600C1808180800201880300C0030;
    char_1900khz[12]  <=   128'h03C0600C300C300C00601880300C0060;
    char_1900khz[13]  <=   128'h03C0600C300C300C00401900300C0060;
    char_1900khz[14]  <=   128'h03C0600C300C300C00C01900300C00C0;
    char_1900khz[15]  <=   128'h03C0600C300C300C00801B00300C00C0;
    char_1900khz[16]  <=   128'h03C0701C300C300C01801D803FFC0180;
    char_1900khz[17]  <=   128'h03C0302C300C300C01001D80300C0180;
    char_1900khz[18]  <=   128'h03C0186C300C300C030018C0300C0300;
    char_1900khz[19]  <=   128'h03C00F8C300C300C020018C0300C0300;
    char_1900khz[20]  <=   128'h03C0000C300C300C06001860300C0600;
    char_1900khz[21]  <=   128'h03C00018300C300C04001860300C0600;
    char_1900khz[22]  <=   128'h03C00018180818080C001830300C0C00;
    char_1900khz[23]  <=   128'h03C000101818181808001830300C1802;
    char_1900khz[24]  <=   128'h03C030301818181818001830300C1806;
    char_1900khz[25]  <=   128'h03C030600C300C3010001818300C3004;
    char_1900khz[26]  <=   128'h03E030C00620062030001818300C301C;
    char_1900khz[27]  <=   128'h1FFC0F8003C003C020007E3EFC3F7FFC;
    char_1900khz[28]  <=   128'h00000000000000006000000000000000;
    char_1900khz[29]  <=   128'h00000000000000004000000000000000;
    char_1900khz[30]  <=   128'h00000000000000000000000000000000;
    char_1900khz[31]  <=   128'h00000000000000000000000000000000;
end 

reg [47:0] char_3d3 [31:0];
                            //空2空 对应MHZ级别
                               always @(posedge lcd_pclk) begin
                                char_3d3[0 ]  <=   48'h000000000000;
                                char_3d3[1 ]  <=   48'h000000000000;
                                char_3d3[2 ]  <=   48'h000000000000;
                                char_3d3[3 ]  <=   48'h000000000000;
                                char_3d3[4 ]  <=   48'h000000000000;
                                char_3d3[5 ]  <=   48'h000000000000;
                                char_3d3[6 ]  <=   48'h07C0000007C0;
                                char_3d3[7 ]  <=   48'h186000001860;
                                char_3d3[8 ]  <=   48'h303000003030;
                                char_3d3[9 ]  <=   48'h301800003018;
                                char_3d3[10]  <=   48'h301800003018;
                                char_3d3[11]  <=   48'h301800003018;
                                char_3d3[12]  <=   48'h001800000018;
                                char_3d3[13]  <=   48'h001800000018;
                                char_3d3[14]  <=   48'h003000000030;
                                char_3d3[15]  <=   48'h006000000060;
                                char_3d3[16]  <=   48'h03C0000003C0;
                                char_3d3[17]  <=   48'h007000000070;
                                char_3d3[18]  <=   48'h001800000018;
                                char_3d3[19]  <=   48'h000800000008;
                                char_3d3[20]  <=   48'h000C0000000C;
                                char_3d3[21]  <=   48'h000C0000000C;
                                char_3d3[22]  <=   48'h300C0000300C;
                                char_3d3[23]  <=   48'h300C0000300C;
                                char_3d3[24]  <=   48'h300818003008;
                                char_3d3[25]  <=   48'h30183C003018;
                                char_3d3[26]  <=   48'h18303C001830;
                                char_3d3[27]  <=   48'h07C0180007C0;
                                char_3d3[28]  <=   48'h000000000000;
                                char_3d3[29]  <=   48'h000000000000;
                                char_3d3[30]  <=   48'h000000000000;
                                char_3d3[31]  <=   48'h000000000000;
                        end 
                            
                        reg [47:0] char_k3k [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_k3k[0 ]  <=   48'h000000000000;
                            char_k3k[1 ]  <=   48'h000000000000;
                            char_k3k[2 ]  <=   48'h000000000000;
                            char_k3k[3 ]  <=   48'h000000000000;
                            char_k3k[4 ]  <=   48'h000000000000;
                            char_k3k[5 ]  <=   48'h000000000000;
                            char_k3k[6 ]  <=   48'h000007C00000;
                            char_k3k[7 ]  <=   48'h000018600000;
                            char_k3k[8 ]  <=   48'h000030300000;
                            char_k3k[9 ]  <=   48'h000030180000;
                            char_k3k[10]  <=   48'h000030180000;
                            char_k3k[11]  <=   48'h000030180000;
                            char_k3k[12]  <=   48'h000000180000;
                            char_k3k[13]  <=   48'h000000180000;
                            char_k3k[14]  <=   48'h000000300000;
                            char_k3k[15]  <=   48'h000000600000;
                            char_k3k[16]  <=   48'h000003C00000;
                            char_k3k[17]  <=   48'h000000700000;
                            char_k3k[18]  <=   48'h000000180000;
                            char_k3k[19]  <=   48'h000000080000;
                            char_k3k[20]  <=   48'h0000000C0000;
                            char_k3k[21]  <=   48'h0000000C0000;
                            char_k3k[22]  <=   48'h0000300C0000;
                            char_k3k[23]  <=   48'h0000300C0000;
                            char_k3k[24]  <=   48'h000030080000;
                            char_k3k[25]  <=   48'h000030180000;
                            char_k3k[26]  <=   48'h000018300000;
                            char_k3k[27]  <=   48'h000007C00000;
                            char_k3k[28]  <=   48'h000000000000;
                            char_k3k[29]  <=   48'h000000000000;
                            char_k3k[30]  <=   48'h000000000000;
                            char_k3k[31]  <=   48'h000000000000;
                        end 
                        
                        
                        reg [47:0] char_k5k [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_k5k[0 ]  <=   48'h000000000000;
                            char_k5k[1 ]  <=   48'h000000000000;
                            char_k5k[2 ]  <=   48'h000000000000;
                            char_k5k[3 ]  <=   48'h000000000000;
                            char_k5k[4 ]  <=   48'h000000000000;
                            char_k5k[5 ]  <=   48'h000000000000;
                            char_k5k[6 ]  <=   48'h00000FFC0000;
                            char_k5k[7 ]  <=   48'h00000FFC0000;
                            char_k5k[8 ]  <=   48'h000010000000;
                            char_k5k[9 ]  <=   48'h000010000000;
                            char_k5k[10]  <=   48'h000010000000;
                            char_k5k[11]  <=   48'h000010000000;
                            char_k5k[12]  <=   48'h000010000000;
                            char_k5k[13]  <=   48'h000010000000;
                            char_k5k[14]  <=   48'h000013E00000;
                            char_k5k[15]  <=   48'h000014300000;
                            char_k5k[16]  <=   48'h000018180000;
                            char_k5k[17]  <=   48'h000010080000;
                            char_k5k[18]  <=   48'h0000000C0000;
                            char_k5k[19]  <=   48'h0000000C0000;
                            char_k5k[20]  <=   48'h0000000C0000;
                            char_k5k[21]  <=   48'h0000000C0000;
                            char_k5k[22]  <=   48'h0000300C0000;
                            char_k5k[23]  <=   48'h0000300C0000;
                            char_k5k[24]  <=   48'h000020180000;
                            char_k5k[25]  <=   48'h000020180000;
                            char_k5k[26]  <=   48'h000018300000;
                            char_k5k[27]  <=   48'h000007C00000;
                            char_k5k[28]  <=   48'h000000000000;
                            char_k5k[29]  <=   48'h000000000000;
                            char_k5k[30]  <=   48'h000000000000;
                            char_k5k[31]  <=   48'h000000000000;
                        end 
                        
                        reg [47:0] char_6d7 [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_6d7[0 ]  <=   48'h000000000000;
                            char_6d7[1 ]  <=   48'h000000000000;
                            char_6d7[2 ]  <=   48'h000000000000;
                            char_6d7[3 ]  <=   48'h000000000000;
                            char_6d7[4 ]  <=   48'h000000000000;
                            char_6d7[5 ]  <=   48'h000000000000;
                            char_6d7[6 ]  <=   48'h01E000001FFC;
                            char_6d7[7 ]  <=   48'h061800001FFC;
                            char_6d7[8 ]  <=   48'h0C1800001008;
                            char_6d7[9 ]  <=   48'h081800003010;
                            char_6d7[10]  <=   48'h180000002010;
                            char_6d7[11]  <=   48'h100000002020;
                            char_6d7[12]  <=   48'h100000000020;
                            char_6d7[13]  <=   48'h300000000040;
                            char_6d7[14]  <=   48'h33E000000040;
                            char_6d7[15]  <=   48'h363000000040;
                            char_6d7[16]  <=   48'h381800000080;
                            char_6d7[17]  <=   48'h380800000080;
                            char_6d7[18]  <=   48'h300C00000100;
                            char_6d7[19]  <=   48'h300C00000100;
                            char_6d7[20]  <=   48'h300C00000100;
                            char_6d7[21]  <=   48'h300C00000100;
                            char_6d7[22]  <=   48'h300C00000300;
                            char_6d7[23]  <=   48'h180C00000300;
                            char_6d7[24]  <=   48'h180818000300;
                            char_6d7[25]  <=   48'h0C183C000300;
                            char_6d7[26]  <=   48'h0E303C000300;
                            char_6d7[27]  <=   48'h03E018000300;
                            char_6d7[28]  <=   48'h000000000000;
                            char_6d7[29]  <=   48'h000000000000;
                            char_6d7[30]  <=   48'h000000000000;
                            char_6d7[31]  <=   48'h000000000000;
                        end 
                        
                        reg [47:0] char_kong10 [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_kong10[0 ]  <=   48'h000000000000;
                            char_kong10[1 ]  <=   48'h000000000000;
                            char_kong10[2 ]  <=   48'h000000000000;
                            char_kong10[3 ]  <=   48'h000000000000;
                            char_kong10[4 ]  <=   48'h000000000000;
                            char_kong10[5 ]  <=   48'h000000000000;
                            char_kong10[6 ]  <=   48'h0000008003C0;
                            char_kong10[7 ]  <=   48'h000001800620;
                            char_kong10[8 ]  <=   48'h00001F800C30;
                            char_kong10[9 ]  <=   48'h000001801818;
                            char_kong10[10]  <=   48'h000001801818;
                            char_kong10[11]  <=   48'h000001801808;
                            char_kong10[12]  <=   48'h00000180300C;
                            char_kong10[13]  <=   48'h00000180300C;
                            char_kong10[14]  <=   48'h00000180300C;
                            char_kong10[15]  <=   48'h00000180300C;
                            char_kong10[16]  <=   48'h00000180300C;
                            char_kong10[17]  <=   48'h00000180300C;
                            char_kong10[18]  <=   48'h00000180300C;
                            char_kong10[19]  <=   48'h00000180300C;
                            char_kong10[20]  <=   48'h00000180300C;
                            char_kong10[21]  <=   48'h00000180300C;
                            char_kong10[22]  <=   48'h000001801808;
                            char_kong10[23]  <=   48'h000001801818;
                            char_kong10[24]  <=   48'h000001801818;
                            char_kong10[25]  <=   48'h000001800C30;
                            char_kong10[26]  <=   48'h000003C00620;
                            char_kong10[27]  <=   48'h00001FF803C0;
                            char_kong10[28]  <=   48'h000000000000;
                            char_kong10[29]  <=   48'h000000000000;
                            char_kong10[30]  <=   48'h000000000000;
                            char_kong10[31]  <=   48'h000000000000;
                        end 
                        
                        
                        
                        
                        reg [111:0] char_7d5k [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_7d5k[0 ]  <=   112'h0000000000000000000000000000;
                            char_7d5k[1 ]  <=   112'h0000000000000000000000000000;
                            char_7d5k[2 ]  <=   112'h0000000000000000000000000000;
                            char_7d5k[3 ]  <=   112'h0000000000000002000000000000;
                            char_7d5k[4 ]  <=   112'h0000000000000006000000000000;
                            char_7d5k[5 ]  <=   112'h0000000000000004000000000000;
                            char_7d5k[6 ]  <=   112'h1FFC00000FFC000C7E7CFC3F1FFE;
                            char_7d5k[7 ]  <=   112'h1FFC00000FFC00081830300C1C0C;
                            char_7d5k[8 ]  <=   112'h10080000100000181820300C180C;
                            char_7d5k[9 ]  <=   112'h30100000100000101860300C3018;
                            char_7d5k[10]  <=   112'h20100000100000301840300C2018;
                            char_7d5k[11]  <=   112'h20200000100000201880300C0030;
                            char_7d5k[12]  <=   112'h00200000100000601880300C0060;
                            char_7d5k[13]  <=   112'h00400000100000401900300C0060;
                            char_7d5k[14]  <=   112'h0040000013E000C01900300C00C0;
                            char_7d5k[15]  <=   112'h00400000143000801B00300C00C0;
                            char_7d5k[16]  <=   112'h00800000181801801D803FFC0180;
                            char_7d5k[17]  <=   112'h00800000100801001D80300C0180;
                            char_7d5k[18]  <=   112'h01000000000C030018C0300C0300;
                            char_7d5k[19]  <=   112'h01000000000C020018C0300C0300;
                            char_7d5k[20]  <=   112'h01000000000C06001860300C0600;
                            char_7d5k[21]  <=   112'h01000000000C04001860300C0600;
                            char_7d5k[22]  <=   112'h03000000300C0C001830300C0C00;
                            char_7d5k[23]  <=   112'h03000000300C08001830300C1802;
                            char_7d5k[24]  <=   112'h03001800201818001830300C1806;
                            char_7d5k[25]  <=   112'h03003C00201810001818300C3004;
                            char_7d5k[26]  <=   112'h03003C00183030001818300C301C;
                            char_7d5k[27]  <=   112'h0300180007C020007E3EFC3F7FFC;
                            char_7d5k[28]  <=   112'h0000000000006000000000000000;
                            char_7d5k[29]  <=   112'h0000000000004000000000000000;
                            char_7d5k[30]  <=   112'h0000000000000000000000000000;
                            char_7d5k[31]  <=   112'h0000000000000000000000000000;
                        end 
                        
                        
                        reg [111:0] char_4d5m [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_4d5m[0 ]  <=   112'h0000000000000000000000000000;
                            char_4d5m[1 ]  <=   112'h0000000000000000000000000000;
                            char_4d5m[2 ]  <=   112'h0000000000000000000000000000;
                            char_4d5m[3 ]  <=   112'h0000000000000002000000000000;
                            char_4d5m[4 ]  <=   112'h0000000000000006000000000000;
                            char_4d5m[5 ]  <=   112'h0000000000000004000000000000;
                            char_4d5m[6 ]  <=   112'h006000000FFC000CF00FFC3F1FFE;
                            char_4d5m[7 ]  <=   112'h006000000FFC0008381C300C1C0C;
                            char_4d5m[8 ]  <=   112'h00E0000010000018381C300C180C;
                            char_4d5m[9 ]  <=   112'h00E0000010000010381C300C3018;
                            char_4d5m[10]  <=   112'h0160000010000030381C300C2018;
                            char_4d5m[11]  <=   112'h0160000010000020382C300C0030;
                            char_4d5m[12]  <=   112'h02600000100000602C2C300C0060;
                            char_4d5m[13]  <=   112'h04600000100000402C2C300C0060;
                            char_4d5m[14]  <=   112'h0460000013E000C02C2C300C00C0;
                            char_4d5m[15]  <=   112'h08600000143000802C4C300C00C0;
                            char_4d5m[16]  <=   112'h08600000181801802C4C3FFC0180;
                            char_4d5m[17]  <=   112'h1060000010080100264C300C0180;
                            char_4d5m[18]  <=   112'h30600000000C0300264C300C0300;
                            char_4d5m[19]  <=   112'h20600000000C0200264C300C0300;
                            char_4d5m[20]  <=   112'h40600000000C0600268C300C0600;
                            char_4d5m[21]  <=   112'h7FFC0000000C0400228C300C0600;
                            char_4d5m[22]  <=   112'h00600000300C0C00238C300C0C00;
                            char_4d5m[23]  <=   112'h00600000300C0800238C300C1802;
                            char_4d5m[24]  <=   112'h0060180020181800230C300C1806;
                            char_4d5m[25]  <=   112'h00603C0020181000230C300C3004;
                            char_4d5m[26]  <=   112'h00603C0018303000210C300C301C;
                            char_4d5m[27]  <=   112'h03FC180007C02000F13FFC3F7FFC;
                            char_4d5m[28]  <=   112'h0000000000006000000000000000;
                            char_4d5m[29]  <=   112'h0000000000004000000000000000;
                            char_4d5m[30]  <=   112'h0000000000000000000000000000;
                            char_4d5m[31]  <=   112'h0000000000000000000000000000;
                        end 
                        
                        
                        reg [111:0] char_10mhz [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_10mhz[0 ]  <=   112'h0000000000000000000000000000;
                            char_10mhz[1 ]  <=   112'h0000000000000000000000000000;
                            char_10mhz[2 ]  <=   112'h0000000000000000000000000000;
                            char_10mhz[3 ]  <=   112'h0000000000000002000000000000;
                            char_10mhz[4 ]  <=   112'h0000000000000006000000000000;
                            char_10mhz[5 ]  <=   112'h0000000000000004000000000000;
                            char_10mhz[6 ]  <=   112'h0000008003C0000CF00FFC3F1FFE;
                            char_10mhz[7 ]  <=   112'h0000018006200008381C300C1C0C;
                            char_10mhz[8 ]  <=   112'h00001F800C300018381C300C180C;
                            char_10mhz[9 ]  <=   112'h0000018018180010381C300C3018;
                            char_10mhz[10]  <=   112'h0000018018180030381C300C2018;
                            char_10mhz[11]  <=   112'h0000018018080020382C300C0030;
                            char_10mhz[12]  <=   112'h00000180300C00602C2C300C0060;
                            char_10mhz[13]  <=   112'h00000180300C00402C2C300C0060;
                            char_10mhz[14]  <=   112'h00000180300C00C02C2C300C00C0;
                            char_10mhz[15]  <=   112'h00000180300C00802C4C300C00C0;
                            char_10mhz[16]  <=   112'h00000180300C01802C4C3FFC0180;
                            char_10mhz[17]  <=   112'h00000180300C0100264C300C0180;
                            char_10mhz[18]  <=   112'h00000180300C0300264C300C0300;
                            char_10mhz[19]  <=   112'h00000180300C0200264C300C0300;
                            char_10mhz[20]  <=   112'h00000180300C0600268C300C0600;
                            char_10mhz[21]  <=   112'h00000180300C0400228C300C0600;
                            char_10mhz[22]  <=   112'h0000018018080C00238C300C0C00;
                            char_10mhz[23]  <=   112'h0000018018180800238C300C1802;
                            char_10mhz[24]  <=   112'h0000018018181800230C300C1806;
                            char_10mhz[25]  <=   112'h000001800C301000230C300C3004;
                            char_10mhz[26]  <=   112'h000003C006203000210C300C301C;
                            char_10mhz[27]  <=   112'h00001FF803C02000F13FFC3F7FFC;
                            char_10mhz[28]  <=   112'h0000000000006000000000000000;
                            char_10mhz[29]  <=   112'h0000000000004000000000000000;
                            char_10mhz[30]  <=   112'h0000000000000000000000000000;
                            char_10mhz[31]  <=   112'h0000000000000000000000000000;
                        end 
                        
                        
                        
                                
                        
                        reg [111:0] char_15khz [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_15khz[0 ]  <=   112'h0000000000000000000000000000;
                            char_15khz[1 ]  <=   112'h0000000000000000000000000000;
                            char_15khz[2 ]  <=   112'h0000000000000000000000000000;
                            char_15khz[3 ]  <=   112'h0000000000000002000000000000;
                            char_15khz[4 ]  <=   112'h0000000000000006000000000000;
                            char_15khz[5 ]  <=   112'h0000000000000004000000000000;
                            char_15khz[6 ]  <=   112'h000000800FFC000C7E7CFC3F1FFE;
                            char_15khz[7 ]  <=   112'h000001800FFC00081830300C1C0C;
                            char_15khz[8 ]  <=   112'h00001F80100000181820300C180C;
                            char_15khz[9 ]  <=   112'h00000180100000101860300C3018;
                            char_15khz[10]  <=   112'h00000180100000301840300C2018;
                            char_15khz[11]  <=   112'h00000180100000201880300C0030;
                            char_15khz[12]  <=   112'h00000180100000601880300C0060;
                            char_15khz[13]  <=   112'h00000180100000401900300C0060;
                            char_15khz[14]  <=   112'h0000018013E000C01900300C00C0;
                            char_15khz[15]  <=   112'h00000180143000801B00300C00C0;
                            char_15khz[16]  <=   112'h00000180181801801D803FFC0180;
                            char_15khz[17]  <=   112'h00000180100801001D80300C0180;
                            char_15khz[18]  <=   112'h00000180000C030018C0300C0300;
                            char_15khz[19]  <=   112'h00000180000C020018C0300C0300;
                            char_15khz[20]  <=   112'h00000180000C06001860300C0600;
                            char_15khz[21]  <=   112'h00000180000C04001860300C0600;
                            char_15khz[22]  <=   112'h00000180300C0C001830300C0C00;
                            char_15khz[23]  <=   112'h00000180300C08001830300C1802;
                            char_15khz[24]  <=   112'h00000180201818001830300C1806;
                            char_15khz[25]  <=   112'h00000180201810001818300C3004;
                            char_15khz[26]  <=   112'h000003C0183030001818300C301C;
                            char_15khz[27]  <=   112'h00001FF807C020007E3EFC3F7FFC;
                            char_15khz[28]  <=   112'h0000000000006000000000000000;
                            char_15khz[29]  <=   112'h0000000000004000000000000000;
                            char_15khz[30]  <=   112'h0000000000000000000000000000;
                            char_15khz[31]  <=   112'h0000000000000000000000000000;
                        end 
                        
                        reg [111:0] char_30khz [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_30khz[0 ]  <=   112'h0000000000000000000000000000;
                            char_30khz[1 ]  <=   112'h0000000000000000000000000000;
                            char_30khz[2 ]  <=   112'h0000000000000000000000000000;
                            char_30khz[3 ]  <=   112'h0000000000000002000000000000;
                            char_30khz[4 ]  <=   112'h0000000000000006000000000000;
                            char_30khz[5 ]  <=   112'h0000000000000004000000000000;
                            char_30khz[6 ]  <=   112'h000007C003C0000C7E7CFC3F1FFE;
                            char_30khz[7 ]  <=   112'h00001860062000081830300C1C0C;
                            char_30khz[8 ]  <=   112'h000030300C3000181820300C180C;
                            char_30khz[9 ]  <=   112'h00003018181800101860300C3018;
                            char_30khz[10]  <=   112'h00003018181800301840300C2018;
                            char_30khz[11]  <=   112'h00003018180800201880300C0030;
                            char_30khz[12]  <=   112'h00000018300C00601880300C0060;
                            char_30khz[13]  <=   112'h00000018300C00401900300C0060;
                            char_30khz[14]  <=   112'h00000030300C00C01900300C00C0;
                            char_30khz[15]  <=   112'h00000060300C00801B00300C00C0;
                            char_30khz[16]  <=   112'h000003C0300C01801D803FFC0180;
                            char_30khz[17]  <=   112'h00000070300C01001D80300C0180;
                            char_30khz[18]  <=   112'h00000018300C030018C0300C0300;
                            char_30khz[19]  <=   112'h00000008300C020018C0300C0300;
                            char_30khz[20]  <=   112'h0000000C300C06001860300C0600;
                            char_30khz[21]  <=   112'h0000000C300C04001860300C0600;
                            char_30khz[22]  <=   112'h0000300C18080C001830300C0C00;
                            char_30khz[23]  <=   112'h0000300C181808001830300C1802;
                            char_30khz[24]  <=   112'h00003008181818001830300C1806;
                            char_30khz[25]  <=   112'h000030180C3010001818300C3004;
                            char_30khz[26]  <=   112'h00001830062030001818300C301C;
                            char_30khz[27]  <=   112'h000007C003C020007E3EFC3F7FFC;
                            char_30khz[28]  <=   112'h0000000000006000000000000000;
                            char_30khz[29]  <=   112'h0000000000004000000000000000;
                            char_30khz[30]  <=   112'h0000000000000000000000000000;
                            char_30khz[31]  <=   112'h0000000000000000000000000000;
                        end 
                        
                        
                        
                        reg [63:0] char_680 [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_680[0 ]  <=   64'h0000000000000000;
                            char_680[1 ]  <=   64'h0000000000000000;
                            char_680[2 ]  <=   64'h0000000000000000;
                            char_680[3 ]  <=   64'h0000000000000000;
                            char_680[4 ]  <=   64'h0000000000000000;
                            char_680[5 ]  <=   64'h0000000000000000;
                            char_680[6 ]  <=   64'h000001E007E003C0;
                            char_680[7 ]  <=   64'h000006180C300620;
                            char_680[8 ]  <=   64'h00000C1818180C30;
                            char_680[9 ]  <=   64'h00000818300C1818;
                            char_680[10]  <=   64'h00001800300C1818;
                            char_680[11]  <=   64'h00001000300C1808;
                            char_680[12]  <=   64'h00001000380C300C;
                            char_680[13]  <=   64'h000030003808300C;
                            char_680[14]  <=   64'h000033E01E18300C;
                            char_680[15]  <=   64'h000036300F20300C;
                            char_680[16]  <=   64'h0000381807C0300C;
                            char_680[17]  <=   64'h0000380818F0300C;
                            char_680[18]  <=   64'h0000300C3078300C;
                            char_680[19]  <=   64'h0000300C3038300C;
                            char_680[20]  <=   64'h0000300C601C300C;
                            char_680[21]  <=   64'h0000300C600C300C;
                            char_680[22]  <=   64'h0000300C600C1808;
                            char_680[23]  <=   64'h0000180C600C1818;
                            char_680[24]  <=   64'h00001808600C1818;
                            char_680[25]  <=   64'h00000C1830180C30;
                            char_680[26]  <=   64'h00000E3018300620;
                            char_680[27]  <=   64'h000003E007C003C0;
                            char_680[28]  <=   64'h0000000000000000;
                            char_680[29]  <=   64'h0000000000000000;
                            char_680[30]  <=   64'h0000000000000000;
                            char_680[31]  <=   64'h0000000000000000;
                        end 
                        
                        
                        reg [63:0] char_1350 [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_1350[0 ]  <=   64'h0000000000000000;
                            char_1350[1 ]  <=   64'h0000000000000000;
                            char_1350[2 ]  <=   64'h0000000000000000;
                            char_1350[3 ]  <=   64'h0000000000000000;
                            char_1350[4 ]  <=   64'h0000000000000000;
                            char_1350[5 ]  <=   64'h0000000000000000;
                            char_1350[6 ]  <=   64'h008007C00FFC03C0;
                            char_1350[7 ]  <=   64'h018018600FFC0620;
                            char_1350[8 ]  <=   64'h1F80303010000C30;
                            char_1350[9 ]  <=   64'h0180301810001818;
                            char_1350[10]  <=   64'h0180301810001818;
                            char_1350[11]  <=   64'h0180301810001808;
                            char_1350[12]  <=   64'h018000181000300C;
                            char_1350[13]  <=   64'h018000181000300C;
                            char_1350[14]  <=   64'h0180003013E0300C;
                            char_1350[15]  <=   64'h018000601430300C;
                            char_1350[16]  <=   64'h018003C01818300C;
                            char_1350[17]  <=   64'h018000701008300C;
                            char_1350[18]  <=   64'h01800018000C300C;
                            char_1350[19]  <=   64'h01800008000C300C;
                            char_1350[20]  <=   64'h0180000C000C300C;
                            char_1350[21]  <=   64'h0180000C000C300C;
                            char_1350[22]  <=   64'h0180300C300C1808;
                            char_1350[23]  <=   64'h0180300C300C1818;
                            char_1350[24]  <=   64'h0180300820181818;
                            char_1350[25]  <=   64'h0180301820180C30;
                            char_1350[26]  <=   64'h03C0183018300620;
                            char_1350[27]  <=   64'h1FF807C007C003C0;
                            char_1350[28]  <=   64'h0000000000000000;
                            char_1350[29]  <=   64'h0000000000000000;
                            char_1350[30]  <=   64'h0000000000000000;
                            char_1350[31]  <=   64'h0000000000000000;
                        end 
                        
                        reg [127:0] char_2000khz [31:0];
                        //空2空 对应MHZ级别
                           always @(posedge lcd_pclk) begin
                            char_2000khz[0 ]  <=   128'h00000000000000000000000000000000;
                            char_2000khz[1 ]  <=   128'h00000000000000000000000000000000;
                            char_2000khz[2 ]  <=   128'h00000000000000000000000000000000;
                            char_2000khz[3 ]  <=   128'h00000000000000000002000000000000;
                            char_2000khz[4 ]  <=   128'h00000000000000000006000000000000;
                            char_2000khz[5 ]  <=   128'h00000000000000000004000000000000;
                            char_2000khz[6 ]  <=   128'h0FF003C003C003C0000C7E7CFC3F1FFE;
                            char_2000khz[7 ]  <=   128'h1E7806200620062000081830300C1C0C;
                            char_2000khz[8 ]  <=   128'h383C0C300C300C3000181820300C180C;
                            char_2000khz[9 ]  <=   128'h381C18181818181800101860300C3018;
                            char_2000khz[10]  <=   128'h781C18181818181800301840300C2018;
                            char_2000khz[11]  <=   128'h781C18081808180800201880300C0030;
                            char_2000khz[12]  <=   128'h7C1C300C300C300C00601880300C0060;
                            char_2000khz[13]  <=   128'h381C300C300C300C00401900300C0060;
                            char_2000khz[14]  <=   128'h003C300C300C300C00C01900300C00C0;
                            char_2000khz[15]  <=   128'h0038300C300C300C00801B00300C00C0;
                            char_2000khz[16]  <=   128'h0070300C300C300C01801D803FFC0180;
                            char_2000khz[17]  <=   128'h00F0300C300C300C01001D80300C0180;
                            char_2000khz[18]  <=   128'h01E0300C300C300C030018C0300C0300;
                            char_2000khz[19]  <=   128'h03C0300C300C300C020018C0300C0300;
                            char_2000khz[20]  <=   128'h0780300C300C300C06001860300C0600;
                            char_2000khz[21]  <=   128'h0F00300C300C300C04001860300C0600;
                            char_2000khz[22]  <=   128'h0E061808180818080C001830300C0C00;
                            char_2000khz[23]  <=   128'h1C0E18181818181808001830300C1802;
                            char_2000khz[24]  <=   128'h380C18181818181818001830300C1806;
                            char_2000khz[25]  <=   128'h701C0C300C300C3010001818300C3004;
                            char_2000khz[26]  <=   128'h7FFC06200620062030001818300C301C;
                            char_2000khz[27]  <=   128'h7FFC03C003C003C020007E3EFC3F7FFC;
                            char_2000khz[28]  <=   128'h00000000000000006000000000000000;
                            char_2000khz[29]  <=   128'h00000000000000004000000000000000;
                            char_2000khz[30]  <=   128'h00000000000000000000000000000000;
                            char_2000khz[31]  <=   128'h00000000000000000000000000000000;
                        end 
                        
                  

reg [47:0] char_2MHZ [31:0];
//空2空 对应MHZ级别
   always @(posedge lcd_pclk) begin
    char_2MHZ[0 ]  <=   48'h000000000000;
    char_2MHZ[1 ]  <=   48'h000000000000;
    char_2MHZ[2 ]  <=   48'h000000000000;
    char_2MHZ[3 ]  <=   48'h000000000000;
    char_2MHZ[4 ]  <=   48'h000000000000;
    char_2MHZ[5 ]  <=   48'h000000000000;
    char_2MHZ[6 ]  <=   48'h000007E00000;
    char_2MHZ[7 ]  <=   48'h000008380000;
    char_2MHZ[8 ]  <=   48'h000010180000;
    char_2MHZ[9 ]  <=   48'h0000200C0000;
    char_2MHZ[10]  <=   48'h0000200C0000;
    char_2MHZ[11]  <=   48'h0000300C0000;
    char_2MHZ[12]  <=   48'h0000300C0000;
    char_2MHZ[13]  <=   48'h0000000C0000;
    char_2MHZ[14]  <=   48'h000000180000;
    char_2MHZ[15]  <=   48'h000000180000;
    char_2MHZ[16]  <=   48'h000000300000;
    char_2MHZ[17]  <=   48'h000000600000;
    char_2MHZ[18]  <=   48'h000000C00000;
    char_2MHZ[19]  <=   48'h000001800000;
    char_2MHZ[20]  <=   48'h000003000000;
    char_2MHZ[21]  <=   48'h000002000000;
    char_2MHZ[22]  <=   48'h000004040000;
    char_2MHZ[23]  <=   48'h000008040000;
    char_2MHZ[24]  <=   48'h000010040000;
    char_2MHZ[25]  <=   48'h0000200C0000;
    char_2MHZ[26]  <=   48'h00003FF80000;
    char_2MHZ[27]  <=   48'h00003FF80000;
    char_2MHZ[28]  <=   48'h000000000000;
    char_2MHZ[29]  <=   48'h000000000000;
    char_2MHZ[30]  <=   48'h000000000000;
    char_2MHZ[31]  <=   48'h000000000000;
    end 


    reg [111:0] char_6MHZ [31:0];
    //空6空 mhz 对应MHZ级别
always @(posedge lcd_pclk) begin
        char_6MHZ[0 ]  <=   112'h0000000000000000000000000000;
        char_6MHZ[1 ]  <=   112'h0000000000000000000000000000;
        char_6MHZ[2 ]  <=   112'h0000000000000000000000000000;
        char_6MHZ[3 ]  <=   112'h0000000000000002000000000000;
        char_6MHZ[4 ]  <=   112'h0000000000000006000000000000;
        char_6MHZ[5 ]  <=   112'h0000000000000004000000000000;
        char_6MHZ[6 ]  <=   112'h000001E00000000CF00FFC3F1FFE;
        char_6MHZ[7 ]  <=   112'h0000061800000008381C300C1C0C;
        char_6MHZ[8 ]  <=   112'h00000C1800000018381C300C180C;
        char_6MHZ[9 ]  <=   112'h0000081800000010381C300C3018;
        char_6MHZ[10]  <=   112'h0000180000000030381C300C2018;
        char_6MHZ[11]  <=   112'h0000100000000020382C300C0030;
        char_6MHZ[12]  <=   112'h00001000000000602C2C300C0060;
        char_6MHZ[13]  <=   112'h00003000000000402C2C300C0060;
        char_6MHZ[14]  <=   112'h000033E0000000C02C2C300C00C0;
        char_6MHZ[15]  <=   112'h00003630000000802C4C300C00C0;
        char_6MHZ[16]  <=   112'h00003818000001802C4C3FFC0180;
        char_6MHZ[17]  <=   112'h0000380800000100264C300C0180;
        char_6MHZ[18]  <=   112'h0000300C00000300264C300C0300;
        char_6MHZ[19]  <=   112'h0000300C00000200264C300C0300;
        char_6MHZ[20]  <=   112'h0000300C00000600268C300C0600;
        char_6MHZ[21]  <=   112'h0000300C00000400228C300C0600;
        char_6MHZ[22]  <=   112'h0000300C00000C00238C300C0C00;
        char_6MHZ[23]  <=   112'h0000180C00000800238C300C1802;
        char_6MHZ[24]  <=   112'h0000180800001800230C300C1806;
        char_6MHZ[25]  <=   112'h00000C1800001000230C300C3004;
        char_6MHZ[26]  <=   112'h00000E3000003000210C300C301C;
        char_6MHZ[27]  <=   112'h000003E000002000F13FFC3F7FFC;
        char_6MHZ[28]  <=   112'h0000000000006000000000000000;
        char_6MHZ[29]  <=   112'h0000000000004000000000000000;
        char_6MHZ[30]  <=   112'h0000000000000000000000000000;
        char_6MHZ[31]  <=   112'h0000000000000000000000000000;
        end 

reg [47:0] char_4MHZ [31:0];
 //空6空 mhz 对应MHZ级别
always @(posedge lcd_pclk) begin
        char_4MHZ[0 ]  <=   48'h000000000000;
        char_4MHZ[1 ]  <=   48'h000000000000;
        char_4MHZ[2 ]  <=   48'h000000000000;
        char_4MHZ[3 ]  <=   48'h000000000000;
        char_4MHZ[4 ]  <=   48'h000000000000;
        char_4MHZ[5 ]  <=   48'h000000000000;
        char_4MHZ[6 ]  <=   48'h000000600000;
        char_4MHZ[7 ]  <=   48'h000000600000;
        char_4MHZ[8 ]  <=   48'h000000E00000;
        char_4MHZ[9 ]  <=   48'h000000E00000;
        char_4MHZ[10]  <=   48'h000001600000;
        char_4MHZ[11]  <=   48'h000001600000;
        char_4MHZ[12]  <=   48'h000002600000;
        char_4MHZ[13]  <=   48'h000004600000;
        char_4MHZ[14]  <=   48'h000004600000;
        char_4MHZ[15]  <=   48'h000008600000;
        char_4MHZ[16]  <=   48'h000008600000;
        char_4MHZ[17]  <=   48'h000010600000;
        char_4MHZ[18]  <=   48'h000030600000;
        char_4MHZ[19]  <=   48'h000020600000;
        char_4MHZ[20]  <=   48'h000040600000;
        char_4MHZ[21]  <=   48'h00007FFC0000;
        char_4MHZ[22]  <=   48'h000000600000;
        char_4MHZ[23]  <=   48'h000000600000;
        char_4MHZ[24]  <=   48'h000000600000;
        char_4MHZ[25]  <=   48'h000000600000;
        char_4MHZ[26]  <=   48'h000000600000;
        char_4MHZ[27]  <=   48'h000003FC0000;
        char_4MHZ[28]  <=   48'h000000000000;
        char_4MHZ[29]  <=   48'h000000000000;
        char_4MHZ[30]  <=   48'h000000000000;
        char_4MHZ[31]  <=   48'h000000000000;
        end 
    
        reg [111:0] char_15MHZ [31:0];
        //空4空 mhz 对应MHZ级别
  always @(posedge lcd_pclk) begin
          char_15MHZ[0 ]  <=   112'h0000000000000000000000000000;
          char_15MHZ[1 ]  <=   112'h0000000000000000000000000000;
          char_15MHZ[2 ]  <=   112'h0000000000000000000000000000;
          char_15MHZ[3 ]  <=   112'h0000000000000002000000000000;
          char_15MHZ[4 ]  <=   112'h0000000000000006000000000000;
          char_15MHZ[5 ]  <=   112'h0000000000000004000000000000;
          char_15MHZ[6 ]  <=   112'h000000800FFC000CF00FFC3F1FFE;
          char_15MHZ[7 ]  <=   112'h000001800FFC0008381C300C1C0C;
          char_15MHZ[8 ]  <=   112'h00001F8010000018381C300C180C;
          char_15MHZ[9 ]  <=   112'h0000018010000010381C300C3018;
          char_15MHZ[10]  <=   112'h0000018010000030381C300C2018;
          char_15MHZ[11]  <=   112'h0000018010000020382C300C0030;
          char_15MHZ[12]  <=   112'h00000180100000602C2C300C0060;
          char_15MHZ[13]  <=   112'h00000180100000402C2C300C0060;
          char_15MHZ[14]  <=   112'h0000018013E000C02C2C300C00C0;
          char_15MHZ[15]  <=   112'h00000180143000802C4C300C00C0;
          char_15MHZ[16]  <=   112'h00000180181801802C4C3FFC0180;
          char_15MHZ[17]  <=   112'h0000018010080100264C300C0180;
          char_15MHZ[18]  <=   112'h00000180000C0300264C300C0300;
          char_15MHZ[19]  <=   112'h00000180000C0200264C300C0300;
          char_15MHZ[20]  <=   112'h00000180000C0600268C300C0600;
          char_15MHZ[21]  <=   112'h00000180000C0400228C300C0600;
          char_15MHZ[22]  <=   112'h00000180300C0C00238C300C0C00;
          char_15MHZ[23]  <=   112'h00000180300C0800238C300C1802;
          char_15MHZ[24]  <=   112'h0000018020181800230C300C1806;
          char_15MHZ[25]  <=   112'h0000018020181000230C300C3004;
          char_15MHZ[26]  <=   112'h000003C018303000210C300C301C;
          char_15MHZ[27]  <=   112'h00001FF807C02000F13FFC3F7FFC;
          char_15MHZ[28]  <=   112'h0000000000006000000000000000;
          char_15MHZ[29]  <=   112'h0000000000004000000000000000;
          char_15MHZ[30]  <=   112'h0000000000000000000000000000;
          char_15MHZ[31]  <=   112'h0000000000000000000000000000;
          end 
           
          reg [47:0] char_5MHZ [31:0];
          //空5空 mhz 对应MHZ级别
 always @(posedge lcd_pclk) begin
         char_5MHZ[0 ]  <=   48'h000000000000;
         char_5MHZ[1 ]  <=   48'h000000000000;
         char_5MHZ[2 ]  <=   48'h000000000000;
         char_5MHZ[3 ]  <=   48'h000000000000;
         char_5MHZ[4 ]  <=   48'h000000000000;
         char_5MHZ[5 ]  <=   48'h000000000000;
         char_5MHZ[6 ]  <=   48'h00000FFC0000;
         char_5MHZ[7 ]  <=   48'h00000FFC0000;
         char_5MHZ[8 ]  <=   48'h000010000000;
         char_5MHZ[9 ]  <=   48'h000010000000;
         char_5MHZ[10]  <=   48'h000010000000;
         char_5MHZ[11]  <=   48'h000010000000;
         char_5MHZ[12]  <=   48'h000010000000;
         char_5MHZ[13]  <=   48'h000010000000;
         char_5MHZ[14]  <=   48'h000013E00000;
         char_5MHZ[15]  <=   48'h000014300000;
         char_5MHZ[16]  <=   48'h000018180000;
         char_5MHZ[17]  <=   48'h000010080000;
         char_5MHZ[18]  <=   48'h0000000C0000;
         char_5MHZ[19]  <=   48'h0000000C0000;
         char_5MHZ[20]  <=   48'h0000000C0000;
         char_5MHZ[21]  <=   48'h0000000C0000;
         char_5MHZ[22]  <=   48'h0000300C0000;
         char_5MHZ[23]  <=   48'h0000300C0000;
         char_5MHZ[24]  <=   48'h000020180000;
         char_5MHZ[25]  <=   48'h000020180000;
         char_5MHZ[26]  <=   48'h000018300000;
         char_5MHZ[27]  <=   48'h000007C00000;
         char_5MHZ[28]  <=   48'h000000000000;
         char_5MHZ[29]  <=   48'h000000000000;
         char_5MHZ[30]  <=   48'h000000000000;
         char_5MHZ[31]  <=   48'h000000000000;
end 

reg [47:0] char_10MHZ [31:0];
//空10  mhz 对应MHZ级别
always @(posedge lcd_pclk) begin
char_10MHZ[0 ]  <=   48'h000000000000;
char_10MHZ[1 ]  <=   48'h000000000000;
char_10MHZ[2 ]  <=   48'h000000000000;
char_10MHZ[3 ]  <=   48'h000000000000;
char_10MHZ[4 ]  <=   48'h000000000000;
char_10MHZ[5 ]  <=   48'h000000000000;
char_10MHZ[6 ]  <=   48'h0000008003C0;
char_10MHZ[7 ]  <=   48'h000001800620;
char_10MHZ[8 ]  <=   48'h00001F800C30;
char_10MHZ[9 ]  <=   48'h000001801818;
char_10MHZ[10]  <=   48'h000001801818;
char_10MHZ[11]  <=   48'h000001801808;
char_10MHZ[12]  <=   48'h00000180300C;
char_10MHZ[13]  <=   48'h00000180300C;
char_10MHZ[14]  <=   48'h00000180300C;
char_10MHZ[15]  <=   48'h00000180300C;
char_10MHZ[16]  <=   48'h00000180300C;
char_10MHZ[17]  <=   48'h00000180300C;
char_10MHZ[18]  <=   48'h00000180300C;
char_10MHZ[19]  <=   48'h00000180300C;
char_10MHZ[20]  <=   48'h00000180300C;
char_10MHZ[21]  <=   48'h00000180300C;
char_10MHZ[22]  <=   48'h000001801808;
char_10MHZ[23]  <=   48'h000001801818;
char_10MHZ[24]  <=   48'h000001801818;
char_10MHZ[25]  <=   48'h000001800C30;
char_10MHZ[26]  <=   48'h000003C00620;
char_10MHZ[27]  <=   48'h00001FF803C0;
char_10MHZ[28]  <=   48'h000000000000;
char_10MHZ[29]  <=   48'h000000000000;
char_10MHZ[30]  <=   48'h000000000000;
char_10MHZ[31]  <=   48'h000000000000;
end 
/*
reg [47:0] char_333 [31:0];
//333   对应KHZ级别
always @(posedge lcd_pclk) begin
char_333[0 ]  <=   48'h000000000000;
char_333[1 ]  <=   48'h000000000000;
char_333[2 ]  <=   48'h000000000000;
char_333[3 ]  <=   48'h000000000000;
char_333[4 ]  <=   48'h000000000000;
char_333[5 ]  <=   48'h000000000000;
char_333[6 ]  <=   48'h07C007C007C0;
char_333[7 ]  <=   48'h186018601860;
char_333[8 ]  <=   48'h303030303030;
char_333[9 ]  <=   48'h301830183018;
char_333[10]  <=   48'h301830183018;
char_333[11]  <=   48'h301830183018;
char_333[12]  <=   48'h001800180018;
char_333[13]  <=   48'h001800180018;
char_333[14]  <=   48'h003000300030;
char_333[15]  <=   48'h006000600060;
char_333[16]  <=   48'h03C003C003C0;
char_333[17]  <=   48'h007000700070;
char_333[18]  <=   48'h001800180018;
char_333[19]  <=   48'h000800080008;
char_333[20]  <=   48'h000C000C000C;
char_333[21]  <=   48'h000C000C000C;
char_333[22]  <=   48'h300C300C300C;
char_333[23]  <=   48'h300C300C300C;
char_333[24]  <=   48'h300830083008;
char_333[25]  <=   48'h301830183018;
char_333[26]  <=   48'h183018301830;
char_333[27]  <=   48'h07C007C007C0;
char_333[28]  <=   48'h000000000000;
char_333[29]  <=   48'h000000000000;
char_333[30]  <=   48'h000000000000;
char_333[31]  <=   48'h000000000000;
end 

reg [47:0] char_667 [31:0];
//667  mhz 对应MHZ级别
always @(posedge lcd_pclk) begin
char_667[0 ]  <=   48'h000000000000;
char_667[1 ]  <=   48'h000000000000;
char_667[2 ]  <=   48'h000000000000;
char_667[3 ]  <=   48'h000000000000;
char_667[4 ]  <=   48'h000000000000;
char_667[5 ]  <=   48'h000000000000;
char_667[6 ]  <=   48'h01E001E01FFC;
char_667[7 ]  <=   48'h061806181FFC;
char_667[8 ]  <=   48'h0C180C181008;
char_667[9 ]  <=   48'h081808183010;
char_667[10]  <=   48'h180018002010;
char_667[11]  <=   48'h100010002020;
char_667[12]  <=   48'h100010000020;
char_667[13]  <=   48'h300030000040;
char_667[14]  <=   48'h33E033E00040;
char_667[15]  <=   48'h363036300040;
char_667[16]  <=   48'h381838180080;
char_667[17]  <=   48'h380838080080;
char_667[18]  <=   48'h300C300C0100;
char_667[19]  <=   48'h300C300C0100;
char_667[20]  <=   48'h300C300C0100;
char_667[21]  <=   48'h300C300C0100;
char_667[22]  <=   48'h300C300C0300;
char_667[23]  <=   48'h180C180C0300;
char_667[24]  <=   48'h180818080300;
char_667[25]  <=   48'h0C180C180300;
char_667[26]  <=   48'h0E300E300300;
char_667[27]  <=   48'h03E003E00300;
char_667[28]  <=   48'h000000000000;
char_667[29]  <=   48'h000000000000;
char_667[30]  <=   48'h000000000000;
char_667[31]  <=   48'h000000000000;
end 
*/
reg [127:0] char_1000 [31:0];
//667  mhz 对应MHZ级别
always @(posedge lcd_pclk) begin
char_1000[0 ]  <=   128'h00000000000000000000000000000000;
char_1000[1 ]  <=   128'h00000000000000000000000000000000;
char_1000[2 ]  <=   128'h00000000000000000000000000000000;
char_1000[3 ]  <=   128'h00000000000000000002000000000000;
char_1000[4 ]  <=   128'h00000000000000000006000000000000;
char_1000[5 ]  <=   128'h00000000000000000004000000000000;
char_1000[6 ]  <=   128'h00C003C003C003C0000C7E7CFC3F1FFE;
char_1000[7 ]  <=   128'h03C006200620062000081830300C1C0C;
char_1000[8 ]  <=   128'h1FC00C300C300C3000181820300C180C;
char_1000[9 ]  <=   128'h03C018181818181800101860300C3018;
char_1000[10]  <=   128'h03C018181818181800301840300C2018;
char_1000[11]  <=   128'h03C018081808180800201880300C0030;
char_1000[12]  <=   128'h03C0300C300C300C00601880300C0060;
char_1000[13]  <=   128'h03C0300C300C300C00401900300C0060;
char_1000[14]  <=   128'h03C0300C300C300C00C01900300C00C0;
char_1000[15]  <=   128'h03C0300C300C300C00801B00300C00C0;
char_1000[16]  <=   128'h03C0300C300C300C01801D803FFC0180;
char_1000[17]  <=   128'h03C0300C300C300C01001D80300C0180;
char_1000[18]  <=   128'h03C0300C300C300C030018C0300C0300;
char_1000[19]  <=   128'h03C0300C300C300C020018C0300C0300;
char_1000[20]  <=   128'h03C0300C300C300C06001860300C0600;
char_1000[21]  <=   128'h03C0300C300C300C04001860300C0600;
char_1000[22]  <=   128'h03C01808180818080C001830300C0C00;
char_1000[23]  <=   128'h03C018181818181808001830300C1802;
char_1000[24]  <=   128'h03C018181818181818001830300C1806;
char_1000[25]  <=   128'h03C00C300C300C3010001818300C3004;
char_1000[26]  <=   128'h03E006200620062030001818300C301C;
char_1000[27]  <=   128'h1FFC03C003C003C020007E3EFC3F7FFC;
char_1000[28]  <=   128'h00000000000000006000000000000000;
char_1000[29]  <=   128'h00000000000000004000000000000000;
char_1000[30]  <=   128'h00000000000000000000000000000000;
char_1000[31]  <=   128'h00000000000000000000000000000000;
end 


reg [111:0] char_60KHZ [31:0];
//60/khz 对应MHZ级别
always @(posedge lcd_pclk) begin
char_60KHZ[0 ]  <=   112'h0000000000000000000000000000;
char_60KHZ[1 ]  <=   112'h0000000000000000000000000000;
char_60KHZ[2 ]  <=   112'h0000000000000000000000000000;
char_60KHZ[3 ]  <=   112'h0000000000000002000000000000;
char_60KHZ[4 ]  <=   112'h0000000000000006000000000000;
char_60KHZ[5 ]  <=   112'h0000000000000004000000000000;
char_60KHZ[6 ]  <=   112'h000001E003C0000C7E7CFC3F1FFE;
char_60KHZ[7 ]  <=   112'h00000618062000081830300C1C0C;
char_60KHZ[8 ]  <=   112'h00000C180C3000181820300C180C;
char_60KHZ[9 ]  <=   112'h00000818181800101860300C3018;
char_60KHZ[10]  <=   112'h00001800181800301840300C2018;
char_60KHZ[11]  <=   112'h00001000180800201880300C0030;
char_60KHZ[12]  <=   112'h00001000300C00601880300C0060;
char_60KHZ[13]  <=   112'h00003000300C00401900300C0060;
char_60KHZ[14]  <=   112'h000033E0300C00C01900300C00C0;
char_60KHZ[15]  <=   112'h00003630300C00801B00300C00C0;
char_60KHZ[16]  <=   112'h00003818300C01801D803FFC0180;
char_60KHZ[17]  <=   112'h00003808300C01001D80300C0180;
char_60KHZ[18]  <=   112'h0000300C300C030018C0300C0300;
char_60KHZ[19]  <=   112'h0000300C300C020018C0300C0300;
char_60KHZ[20]  <=   112'h0000300C300C06001860300C0600;
char_60KHZ[21]  <=   112'h0000300C300C04001860300C0600;
char_60KHZ[22]  <=   112'h0000300C18080C001830300C0C00;
char_60KHZ[23]  <=   112'h0000180C181808001830300C1802;
char_60KHZ[24]  <=   112'h00001808181818001830300C1806;
char_60KHZ[25]  <=   112'h00000C180C3010001818300C3004;
char_60KHZ[26]  <=   112'h00000E30062030001818300C301C;
char_60KHZ[27]  <=   112'h000003E003C020007E3EFC3F7FFC;
char_60KHZ[28]  <=   112'h0000000000006000000000000000;
char_60KHZ[29]  <=   112'h0000000000004000000000000000;
char_60KHZ[30]  <=   112'h0000000000000000000000000000;
char_60KHZ[31]  <=   112'h0000000000000000000000000000;
end 


reg [111:0] char_120KHZ [31:0];
//120/khz 对应MHZ级别
always @(posedge lcd_pclk) begin
char_120KHZ[0 ]  <=   112'h0000000000000000000000000000;
char_120KHZ[1 ]  <=   112'h0000000000000000000000000000;
char_120KHZ[2 ]  <=   112'h0000000000000000000000000000;
char_120KHZ[3 ]  <=   112'h0000000000000002000000000000;
char_120KHZ[4 ]  <=   112'h0000000000000006000000000000;
char_120KHZ[5 ]  <=   112'h0000000000000004000000000000;
char_120KHZ[6 ]  <=   112'h008007E003C0000C7E7CFC3F1FFE;
char_120KHZ[7 ]  <=   112'h01800838062000081830300C1C0C;
char_120KHZ[8 ]  <=   112'h1F8010180C3000181820300C180C;
char_120KHZ[9 ]  <=   112'h0180200C181800101860300C3018;
char_120KHZ[10]  <=   112'h0180200C181800301840300C2018;
char_120KHZ[11]  <=   112'h0180300C180800201880300C0030;
char_120KHZ[12]  <=   112'h0180300C300C00601880300C0060;
char_120KHZ[13]  <=   112'h0180000C300C00401900300C0060;
char_120KHZ[14]  <=   112'h01800018300C00C01900300C00C0;
char_120KHZ[15]  <=   112'h01800018300C00801B00300C00C0;
char_120KHZ[16]  <=   112'h01800030300C01801D803FFC0180;
char_120KHZ[17]  <=   112'h01800060300C01001D80300C0180;
char_120KHZ[18]  <=   112'h018000C0300C030018C0300C0300;
char_120KHZ[19]  <=   112'h01800180300C020018C0300C0300;
char_120KHZ[20]  <=   112'h01800300300C06001860300C0600;
char_120KHZ[21]  <=   112'h01800200300C04001860300C0600;
char_120KHZ[22]  <=   112'h0180040418080C001830300C0C00;
char_120KHZ[23]  <=   112'h01800804181808001830300C1802;
char_120KHZ[24]  <=   112'h01801004181818001830300C1806;
char_120KHZ[25]  <=   112'h0180200C0C3010001818300C3004;
char_120KHZ[26]  <=   112'h03C03FF8062030001818300C301C;
char_120KHZ[27]  <=   112'h1FF83FF803C020007E3EFC3F7FFC;
char_120KHZ[28]  <=   112'h0000000000006000000000000000;
char_120KHZ[29]  <=   112'h0000000000004000000000000000;
char_120KHZ[30]  <=   112'h0000000000000000000000000000;
char_120KHZ[31]  <=   112'h0000000000000000000000000000;
end 

reg [111:0] char_240KHZ [31:0];
//120/khz 对应MHZ级别
always @(posedge lcd_pclk) begin
char_240KHZ[0 ]  <=   112'h0000000000000000000000000000;
char_240KHZ[1 ]  <=   112'h0000000000000000000000000000;
char_240KHZ[2 ]  <=   112'h0000000000000000000000000000;
char_240KHZ[3 ]  <=   112'h0000000000000002000000000000;
char_240KHZ[4 ]  <=   112'h0000000000000006000000000000;
char_240KHZ[5 ]  <=   112'h0000000000000004000000000000;
char_240KHZ[6 ]  <=   112'h07E0006003C0000C7E7CFC3F1FFE;
char_240KHZ[7 ]  <=   112'h08380060062000081830300C1C0C;
char_240KHZ[8 ]  <=   112'h101800E00C3000181820300C180C;
char_240KHZ[9 ]  <=   112'h200C00E0181800101860300C3018;
char_240KHZ[10]  <=   112'h200C0160181800301840300C2018;
char_240KHZ[11]  <=   112'h300C0160180800201880300C0030;
char_240KHZ[12]  <=   112'h300C0260300C00601880300C0060;
char_240KHZ[13]  <=   112'h000C0460300C00401900300C0060;
char_240KHZ[14]  <=   112'h00180460300C00C01900300C00C0;
char_240KHZ[15]  <=   112'h00180860300C00801B00300C00C0;
char_240KHZ[16]  <=   112'h00300860300C01801D803FFC0180;
char_240KHZ[17]  <=   112'h00601060300C01001D80300C0180;
char_240KHZ[18]  <=   112'h00C03060300C030018C0300C0300;
char_240KHZ[19]  <=   112'h01802060300C020018C0300C0300;
char_240KHZ[20]  <=   112'h03004060300C06001860300C0600;
char_240KHZ[21]  <=   112'h02007FFC300C04001860300C0600;
char_240KHZ[22]  <=   112'h0404006018080C001830300C0C00;
char_240KHZ[23]  <=   112'h08040060181808001830300C1802;
char_240KHZ[24]  <=   112'h10040060181818001830300C1806;
char_240KHZ[25]  <=   112'h200C00600C3010001818300C3004;
char_240KHZ[26]  <=   112'h3FF80060062030001818300C301C;
char_240KHZ[27]  <=   112'h3FF803FC03C020007E3EFC3F7FFC;
char_240KHZ[28]  <=   112'h0000000000006000000000000000;
char_240KHZ[29]  <=   112'h0000000000004000000000000000;
char_240KHZ[30]  <=   112'h0000000000000000000000000000;
char_240KHZ[31]  <=   112'h0000000000000000000000000000;
end 

reg [111:0] char_480KHZ [31:0];
//120/khz 对应MHZ级别
always @(posedge lcd_pclk) begin
char_480KHZ[0 ]  <=   112'h0000000000000000000000000000;
char_480KHZ[1 ]  <=   112'h0000000000000000000000000000;
char_480KHZ[2 ]  <=   112'h0000000000000000000000000000;
char_480KHZ[3 ]  <=   112'h0000000000000002000000000000;
char_480KHZ[4 ]  <=   112'h0000000000000006000000000000;
char_480KHZ[5 ]  <=   112'h0000000000000004000000000000;
char_480KHZ[6 ]  <=   112'h006007E003C0000C7E7CFC3F1FFE;
char_480KHZ[7 ]  <=   112'h00600C30062000081830300C1C0C;
char_480KHZ[8 ]  <=   112'h00E018180C3000181820300C180C;
char_480KHZ[9 ]  <=   112'h00E0300C181800101860300C3018;
char_480KHZ[10]  <=   112'h0160300C181800301840300C2018;
char_480KHZ[11]  <=   112'h0160300C180800201880300C0030;
char_480KHZ[12]  <=   112'h0260380C300C00601880300C0060;
char_480KHZ[13]  <=   112'h04603808300C00401900300C0060;
char_480KHZ[14]  <=   112'h04601E18300C00C01900300C00C0;
char_480KHZ[15]  <=   112'h08600F20300C00801B00300C00C0;
char_480KHZ[16]  <=   112'h086007C0300C01801D803FFC0180;
char_480KHZ[17]  <=   112'h106018F0300C01001D80300C0180;
char_480KHZ[18]  <=   112'h30603078300C030018C0300C0300;
char_480KHZ[19]  <=   112'h20603038300C020018C0300C0300;
char_480KHZ[20]  <=   112'h4060601C300C06001860300C0600;
char_480KHZ[21]  <=   112'h7FFC600C300C04001860300C0600;
char_480KHZ[22]  <=   112'h0060600C18080C001830300C0C00;
char_480KHZ[23]  <=   112'h0060600C181808001830300C1802;
char_480KHZ[24]  <=   112'h0060600C181818001830300C1806;
char_480KHZ[25]  <=   112'h006030180C3010001818300C3004;
char_480KHZ[26]  <=   112'h00601830062030001818300C301C;
char_480KHZ[27]  <=   112'h03FC07C003C020007E3EFC3F7FFC;
char_480KHZ[28]  <=   112'h0000000000006000000000000000;
char_480KHZ[29]  <=   112'h0000000000004000000000000000;
char_480KHZ[30]  <=   112'h0000000000000000000000000000;
char_480KHZ[31]  <=   112'h0000000000000000000000000000;
end 

reg [47:0] char_160 [31:0];
//160 对应MHZ级别
always @(posedge lcd_pclk) begin
char_160[0 ]  <=   48'h000000000000;
char_160[1 ]  <=   48'h000000000000;
char_160[2 ]  <=   48'h000000000000;
char_160[3 ]  <=   48'h000000000000;
char_160[4 ]  <=   48'h000000000000;
char_160[5 ]  <=   48'h000000000000;
char_160[6 ]  <=   48'h008001E003C0;
char_160[7 ]  <=   48'h018006180620;
char_160[8 ]  <=   48'h1F800C180C30;
char_160[9 ]  <=   48'h018008181818;
char_160[10]  <=   48'h018018001818;
char_160[11]  <=   48'h018010001808;
char_160[12]  <=   48'h01801000300C;
char_160[13]  <=   48'h01803000300C;
char_160[14]  <=   48'h018033E0300C;
char_160[15]  <=   48'h01803630300C;
char_160[16]  <=   48'h01803818300C;
char_160[17]  <=   48'h01803808300C;
char_160[18]  <=   48'h0180300C300C;
char_160[19]  <=   48'h0180300C300C;
char_160[20]  <=   48'h0180300C300C;
char_160[21]  <=   48'h0180300C300C;
char_160[22]  <=   48'h0180300C1808;
char_160[23]  <=   48'h0180180C1818;
char_160[24]  <=   48'h018018081818;
char_160[25]  <=   48'h01800C180C30;
char_160[26]  <=   48'h03C00E300620;
char_160[27]  <=   48'h1FF803E003C0;
char_160[28]  <=   48'h000000000000;
char_160[29]  <=   48'h000000000000;
char_160[30]  <=   48'h000000000000;
char_160[31]  <=   48'h000000000000;
end 


reg [47:0] char_320 [31:0];
//320 对应MHZ级别
always @(posedge lcd_pclk) begin
char_320[0 ]  <=   48'h000000000000;
char_320[1 ]  <=   48'h000000000000;
char_320[2 ]  <=   48'h000000000000;
char_320[3 ]  <=   48'h000000000000;
char_320[4 ]  <=   48'h000000000000;
char_320[5 ]  <=   48'h000000000000;
char_320[6 ]  <=   48'h07C007E003C0;
char_320[7 ]  <=   48'h186008380620;
char_320[8 ]  <=   48'h303010180C30;
char_320[9 ]  <=   48'h3018200C1818;
char_320[10]  <=   48'h3018200C1818;
char_320[11]  <=   48'h3018300C1808;
char_320[12]  <=   48'h0018300C300C;
char_320[13]  <=   48'h0018000C300C;
char_320[14]  <=   48'h00300018300C;
char_320[15]  <=   48'h00600018300C;
char_320[16]  <=   48'h03C00030300C;
char_320[17]  <=   48'h00700060300C;
char_320[18]  <=   48'h001800C0300C;
char_320[19]  <=   48'h00080180300C;
char_320[20]  <=   48'h000C0300300C;
char_320[21]  <=   48'h000C0200300C;
char_320[22]  <=   48'h300C04041808;
char_320[23]  <=   48'h300C08041818;
char_320[24]  <=   48'h300810041818;
char_320[25]  <=   48'h3018200C0C30;
char_320[26]  <=   48'h18303FF80620;
char_320[27]  <=   48'h07C03FF803C0;
char_320[28]  <=   48'h000000000000;
char_320[29]  <=   48'h000000000000;
char_320[30]  <=   48'h000000000000;
char_320[31]  <=   48'h000000000000;
end 

reg [47:0] char_kong20 [31:0];
//kong20 对应MHZ级别
always @(posedge lcd_pclk) begin
char_kong20[0 ]  <=   48'h000000000000;
char_kong20[1 ]  <=   48'h000000000000;
char_kong20[2 ]  <=   48'h000000000000;
char_kong20[3 ]  <=   48'h000000000000;
char_kong20[4 ]  <=   48'h000000000000;
char_kong20[5 ]  <=   48'h000000000000;
char_kong20[6 ]  <=   48'h000007E003C0;
char_kong20[7 ]  <=   48'h000008380620;
char_kong20[8 ]  <=   48'h000010180C30;
char_kong20[9 ]  <=   48'h0000200C1818;
char_kong20[10]  <=   48'h0000200C1818;
char_kong20[11]  <=   48'h0000300C1808;
char_kong20[12]  <=   48'h0000300C300C;
char_kong20[13]  <=   48'h0000000C300C;
char_kong20[14]  <=   48'h00000018300C;
char_kong20[15]  <=   48'h00000018300C;
char_kong20[16]  <=   48'h00000030300C;
char_kong20[17]  <=   48'h00000060300C;
char_kong20[18]  <=   48'h000000C0300C;
char_kong20[19]  <=   48'h00000180300C;
char_kong20[20]  <=   48'h00000300300C;
char_kong20[21]  <=   48'h00000200300C;
char_kong20[22]  <=   48'h000004041808;
char_kong20[23]  <=   48'h000008041818;
char_kong20[24]  <=   48'h000010041818;
char_kong20[25]  <=   48'h0000200C0C30;
char_kong20[26]  <=   48'h00003FF80620;
char_kong20[27]  <=   48'h00003FF803C0;
char_kong20[28]  <=   48'h000000000000;
char_kong20[29]  <=   48'h000000000000;
char_kong20[30]  <=   48'h000000000000;
char_kong20[31]  <=   48'h000000000000;
end 


reg [47:0] char_kong40  [31:0];
//kong40  对应MHZ级别
always @(posedge lcd_pclk) begin
char_kong40[0 ]  <=   48'h000000000000;
char_kong40[1 ]  <=   48'h000000000000;
char_kong40[2 ]  <=   48'h000000000000;
char_kong40[3 ]  <=   48'h000000000000;
char_kong40[4 ]  <=   48'h000000000000;
char_kong40[5 ]  <=   48'h000000000000;
char_kong40[6 ]  <=   48'h0000006003C0;
char_kong40[7 ]  <=   48'h000000600620;
char_kong40[8 ]  <=   48'h000000E00C30;
char_kong40[9 ]  <=   48'h000000E01818;
char_kong40[10]  <=   48'h000001601818;
char_kong40[11]  <=   48'h000001601808;
char_kong40[12]  <=   48'h00000260300C;
char_kong40[13]  <=   48'h00000460300C;
char_kong40[14]  <=   48'h00000460300C;
char_kong40[15]  <=   48'h00000860300C;
char_kong40[16]  <=   48'h00000860300C;
char_kong40[17]  <=   48'h00001060300C;
char_kong40[18]  <=   48'h00003060300C;
char_kong40[19]  <=   48'h00002060300C;
char_kong40[20]  <=   48'h00004060300C;
char_kong40[21]  <=   48'h00007FFC300C;
char_kong40[22]  <=   48'h000000601808;
char_kong40[23]  <=   48'h000000601818;
char_kong40[24]  <=   48'h000000601818;
char_kong40[25]  <=   48'h000000600C30;
char_kong40[26]  <=   48'h000000600620;
char_kong40[27]  <=   48'h000003FC03C0;
char_kong40[28]  <=   48'h000000000000;
char_kong40[29]  <=   48'h000000000000;
char_kong40[30]  <=   48'h000000000000;
char_kong40[31]  <=   48'h000000000000;
end 

reg [47:0] char_kong80  [31:0];
//kong80  对应MHZ级别
always @(posedge lcd_pclk) begin
char_kong80[0 ]  <=   48'h000000000000;
char_kong80[1 ]  <=   48'h000000000000;
char_kong80[2 ]  <=   48'h000000000000;
char_kong80[3 ]  <=   48'h000000000000;
char_kong80[4 ]  <=   48'h000000000000;
char_kong80[5 ]  <=   48'h000000000000;
char_kong80[6 ]  <=   48'h000007E003C0;
char_kong80[7 ]  <=   48'h00000C300620;
char_kong80[8 ]  <=   48'h000018180C30;
char_kong80[9 ]  <=   48'h0000300C1818;
char_kong80[10]  <=   48'h0000300C1818;
char_kong80[11]  <=   48'h0000300C1808;
char_kong80[12]  <=   48'h0000380C300C;
char_kong80[13]  <=   48'h00003808300C;
char_kong80[14]  <=   48'h00001E18300C;
char_kong80[15]  <=   48'h00000F20300C;
char_kong80[16]  <=   48'h000007C0300C;
char_kong80[17]  <=   48'h000018F0300C;
char_kong80[18]  <=   48'h00003078300C;
char_kong80[19]  <=   48'h00003038300C;
char_kong80[20]  <=   48'h0000601C300C;
char_kong80[21]  <=   48'h0000600C300C;
char_kong80[22]  <=   48'h0000600C1808;
char_kong80[23]  <=   48'h0000600C1818;
char_kong80[24]  <=   48'h0000600C1818;
char_kong80[25]  <=   48'h000030180C30;
char_kong80[26]  <=   48'h000018300620;
char_kong80[27]  <=   48'h000007C003C0;
char_kong80[28]  <=   48'h000000000000;
char_kong80[29]  <=   48'h000000000000;
char_kong80[30]  <=   48'h000000000000;
char_kong80[31]  <=   48'h000000000000;
end 

reg [111:0] char_30mhz  [31:0];
//kong80  对应MHZ级别
always @(posedge lcd_pclk) begin
char_30mhz[0 ]  <=   112'h0000000000000000000000000000;
char_30mhz[1 ]  <=   112'h0000000000000000000000000000;
char_30mhz[2 ]  <=   112'h0000000000000000000000000000;
char_30mhz[3 ]  <=   112'h0000000000000002000000000000;
char_30mhz[4 ]  <=   112'h0000000000000006000000000000;
char_30mhz[5 ]  <=   112'h0000000000000004000000000000;
char_30mhz[6 ]  <=   112'h000007C003C0000CF00FFC3F1FFE;
char_30mhz[7 ]  <=   112'h0000186006200008381C300C1C0C;
char_30mhz[8 ]  <=   112'h000030300C300018381C300C180C;
char_30mhz[9 ]  <=   112'h0000301818180010381C300C3018;
char_30mhz[10]  <=   112'h0000301818180030381C300C2018;
char_30mhz[11]  <=   112'h0000301818080020382C300C0030;
char_30mhz[12]  <=   112'h00000018300C00602C2C300C0060;
char_30mhz[13]  <=   112'h00000018300C00402C2C300C0060;
char_30mhz[14]  <=   112'h00000030300C00C02C2C300C00C0;
char_30mhz[15]  <=   112'h00000060300C00802C4C300C00C0;
char_30mhz[16]  <=   112'h000003C0300C01802C4C3FFC0180;
char_30mhz[17]  <=   112'h00000070300C0100264C300C0180;
char_30mhz[18]  <=   112'h00000018300C0300264C300C0300;
char_30mhz[19]  <=   112'h00000008300C0200264C300C0300;
char_30mhz[20]  <=   112'h0000000C300C0600268C300C0600;
char_30mhz[21]  <=   112'h0000000C300C0400228C300C0600;
char_30mhz[22]  <=   112'h0000300C18080C00238C300C0C00;
char_30mhz[23]  <=   112'h0000300C18180800238C300C1802;
char_30mhz[24]  <=   112'h0000300818181800230C300C1806;
char_30mhz[25]  <=   112'h000030180C301000230C300C3004;
char_30mhz[26]  <=   112'h0000183006203000210C300C301C;
char_30mhz[27]  <=   112'h000007C003C02000F13FFC3F7FFC;
char_30mhz[28]  <=   112'h0000000000006000000000000000;
char_30mhz[29]  <=   112'h0000000000004000000000000000;
char_30mhz[30]  <=   112'h0000000000000000000000000000;
char_30mhz[31]  <=   112'h0000000000000000000000000000;
end 

reg [63:0] char_k630  [31:0];
//kong80  对应MHZ级别
always @(posedge lcd_pclk) begin
char_k630[0 ]  <=   64'h0000000000000000;
char_k630[1 ]  <=   64'h0000000000000000;
char_k630[2 ]  <=   64'h0000000000000000;
char_k630[3 ]  <=   64'h0000000000000000;
char_k630[4 ]  <=   64'h0000000000000000;
char_k630[5 ]  <=   64'h0000000000000000;
char_k630[6 ]  <=   64'h000001E007C003C0;
char_k630[7 ]  <=   64'h0000061818600620;
char_k630[8 ]  <=   64'h00000C1830300C30;
char_k630[9 ]  <=   64'h0000081830181818;
char_k630[10]  <=   64'h0000180030181818;
char_k630[11]  <=   64'h0000100030181808;
char_k630[12]  <=   64'h000010000018300C;
char_k630[13]  <=   64'h000030000018300C;
char_k630[14]  <=   64'h000033E00030300C;
char_k630[15]  <=   64'h000036300060300C;
char_k630[16]  <=   64'h0000381803C0300C;
char_k630[17]  <=   64'h000038080070300C;
char_k630[18]  <=   64'h0000300C0018300C;
char_k630[19]  <=   64'h0000300C0008300C;
char_k630[20]  <=   64'h0000300C000C300C;
char_k630[21]  <=   64'h0000300C000C300C;
char_k630[22]  <=   64'h0000300C300C1808;
char_k630[23]  <=   64'h0000180C300C1818;
char_k630[24]  <=   64'h0000180830081818;
char_k630[25]  <=   64'h00000C1830180C30;
char_k630[26]  <=   64'h00000E3018300620;
char_k630[27]  <=   64'h000003E007C003C0;
char_k630[28]  <=   64'h0000000000000000;
char_k630[29]  <=   64'h0000000000000000;
char_k630[30]  <=   64'h0000000000000000;
char_k630[31]  <=   64'h0000000000000000;
end 





always @(posedge lcd_pclk or negedge sys_rst_n ) begin
	if (!sys_rst_n )
		pixel_data <= BACK_COLOR;
	else   
	case(freq_adj)
        12'd4095:    
			if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
			&& (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
				if(char_kong10[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
 					pixel_data <= CHAR_COLOR;    //显示字符 20
				else
					pixel_data <= BACK_COLOR;    //显示字符区域的背景色
			end
			else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
			&& (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
				if(char_kong20[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
					pixel_data <= CHAR_COLOR;    //显示字符 40
				else
					pixel_data <= BACK_COLOR;    //显示字符区域的背景色
			end
			else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
			&& (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
				if(char_30khz[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
					pixel_data <= CHAR_COLOR;    //显示字符 60/KHZ
				else
					pixel_data <= BACK_COLOR;    //显示字符区域的背景色
				end
			else 
				pixel_data <= BACK_COLOR;
			12'd2047:    
			if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
			&& (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
				if(char_k5k[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
                         pixel_data <= CHAR_COLOR;    //显示字符 20
           else
                         pixel_data <= BACK_COLOR;    //显示字符区域的背景色
      end
           else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
              && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                      if(char_kong10[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                         pixel_data <= CHAR_COLOR;    //显示字符 40
           else
                         pixel_data <= BACK_COLOR;    //显示字符区域的背景色
      end
           else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
              && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                      if(char_15khz[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                         pixel_data <= CHAR_COLOR;    //显示字符 60/KHZ
           else
                         pixel_data <= BACK_COLOR;    //显示字符区域的背景色
      end
          else 
              pixel_data <= BACK_COLOR;
              12'd1023:    
              if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
                               && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
                         if(char_kong10[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
                            pixel_data <= CHAR_COLOR;    //显示字符 20
              else
                            pixel_data <= BACK_COLOR;    //显示字符区域的背景色
         end
              else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
                 && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                         if(char_kong20[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                            pixel_data <= CHAR_COLOR;    //显示字符 40
              else
                            pixel_data <= BACK_COLOR;    //显示字符区域的背景色
         end
              else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
                 && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                         if(char_30khz[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                            pixel_data <= CHAR_COLOR;    //显示字符 60/KHZ
              else
                            pixel_data <= BACK_COLOR;    //显示字符区域的背景色
         end
             else 
                 pixel_data <= BACK_COLOR;

    12'd511:    
     if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
                      && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
                if(char_kong20[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
                   pixel_data <= CHAR_COLOR;    //显示字符 20
     else
                   pixel_data <= BACK_COLOR;    //显示字符区域的背景色
end
     else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                if(char_kong40[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                   pixel_data <= CHAR_COLOR;    //显示字符 40
     else
                   pixel_data <= BACK_COLOR;    //显示字符区域的背景色
end
     else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                if(char_60KHZ[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                   pixel_data <= CHAR_COLOR;    //显示字符 60/KHZ
     else
                   pixel_data <= BACK_COLOR;    //显示字符区域的背景色
end
    else 
        pixel_data <= BACK_COLOR;
    
    12'd255:    
    if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
        && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
  if(char_kong40[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
     pixel_data <= CHAR_COLOR;    //显示字符 40
    else
     pixel_data <= BACK_COLOR;    //显示字符区域的背景色
end
    else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
&& (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                  if(char_kong80[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                       pixel_data <= CHAR_COLOR;    //显示字符 80
    else
                       pixel_data <= BACK_COLOR;    //显示字符区域的背景色
end
else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
&& (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                  if(char_120KHZ[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                      pixel_data <= CHAR_COLOR;    //显示字符 60/KHZ
else
                     pixel_data <= BACK_COLOR;    //显示字符区域的背景色
end
else 
                     pixel_data <= BACK_COLOR;
    
                     12'd127:   
                        if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
                                         && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
                                   if(char_kong80[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
                                      pixel_data <= CHAR_COLOR;    //显示字符80
                        else
                                      pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                   end
                        else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
                           && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                                   if(char_160[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                                      pixel_data <= CHAR_COLOR;    //显示字符 160
                        else
                                      pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                   end
                        else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
                           && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                                   if(char_240KHZ[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                                      pixel_data <= CHAR_COLOR;    //显示字符 240/KHZ
                        else
                                      pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                   end
                   else 
                     pixel_data <= BACK_COLOR;
                   12'd63:    
                    if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
                                     && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
                               if(char_160[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
                                  pixel_data <= CHAR_COLOR;    //显示字符 160
                    else
                                  pixel_data <= BACK_COLOR;    //显示字符区域的背景色
               end
                    else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
                       && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                               if(char_320[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                                  pixel_data <= CHAR_COLOR;    //显示字符 320
                    else
                                  pixel_data <= BACK_COLOR;    //显示字符区域的背景色
               end
                    else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
                       && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                               if(char_480KHZ[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                                  pixel_data <= CHAR_COLOR;    //显示字符 480/KHZ
                    else
                                  pixel_data <= BACK_COLOR;    //显示字符区域的背景色
               end
                   else 
                               pixel_data <= BACK_COLOR;
                    12'd31:   
                        if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
                                         && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
                                   if(char_320[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
                                      pixel_data <= CHAR_COLOR;    //显示字符 160
                        else
                                      pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                   end
                        else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
                           && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                                   if(char_640[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                                      pixel_data <= CHAR_COLOR;    //显示字符 320
                        else
                                      pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                   end
                        else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
                           && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                                   if(char_960khz[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                                      pixel_data <= CHAR_COLOR;    //显示字符 1000KHZ
                        else
                                      pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                   end
                        else 
                                       pixel_data <= BACK_COLOR;
                    12'd15:   
                                       if((pixel_xpos >= CHAR_X_START_680 - 1'b1) && (pixel_xpos < CHAR_X_START_680 + CHAR_WIDTH_680 - 1'b1)
                                                        && (pixel_ypos >= CHAR_Y_START_680) && (pixel_ypos < CHAR_Y_START_680 + CHAR_HEIGHT)) begin
                                                  if(char_k630[y_cnt_680][CHAR_WIDTH_680 -1'b1 - x_cnt_680])
                                                     pixel_data <= CHAR_COLOR;    //显示字符 160
                                       else
                                                     pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                                  end
                                       else if((pixel_xpos >= CHAR_X_START_135 - 1'b1) && (pixel_xpos < CHAR_X_START_135 + CHAR_WIDTH_135 - 1'b1)
                                          && (pixel_ypos >= CHAR_Y_START_135) && (pixel_ypos < CHAR_Y_START_135 + CHAR_HEIGHT)) begin
                                                  if(char_1270[y_cnt_135][CHAR_WIDTH_135 -1'b1 - x_cnt_135])
                                                     pixel_data <= CHAR_COLOR;    //显示字符 320
                                       else
                                                     pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                                  end
                                       else if((pixel_xpos >= CHAR_X_START_1000 - 1'b1) && (pixel_xpos < CHAR_X_START_1000 + CHAR_WIDTH_1000 - 1'b1)
                                          && (pixel_ypos >= CHAR_Y_START_1000) && (pixel_ypos < CHAR_Y_START_1000 + CHAR_HEIGHT)) begin
                                                  if(char_1900khz[y_cnt_1000][CHAR_WIDTH_1000 -1'b1 - x_cnt_1000])
                                                     pixel_data <= CHAR_COLOR;    //显示字符 1000KHZ
                                       else
                                                     pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                                  end
                                       else 
                                                      pixel_data <= BACK_COLOR;
                     12'd7:    
                    if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
                                     && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
                               if(char_1d3[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
                                  pixel_data <= CHAR_COLOR;    //显示字符2
                    else
                                  pixel_data <= BACK_COLOR;    //显示字符区域的背景色
               end
                    else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
                       && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                               if(char_2d5[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                                  pixel_data <= CHAR_COLOR;    //显示字符 4
                    else
                                  pixel_data <= BACK_COLOR;    //显示字符区域的背景色
               end
                    else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
                       && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                               if(char_3d8mhz[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                                  pixel_data <= CHAR_COLOR;    //显示字符 6m
                    else
                                  pixel_data <= BACK_COLOR;    //显示字符区域的背景色
               end
                    else 
                                pixel_data <= BACK_COLOR;
           
               12'd3:    
                if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
                                 && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
                           if(char_2d5[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
                              pixel_data <= CHAR_COLOR;    //显示字符 160
                else
                              pixel_data <= BACK_COLOR;    //显示字符区域的背景色
           end
                else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
                   && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                           if(char_k5k[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                              pixel_data <= CHAR_COLOR;    //显示字符 320
                else
                              pixel_data <= BACK_COLOR;    //显示字符区域的背景色
           end
                else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
                   && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                           if(char_7d6mhz[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                              pixel_data <= CHAR_COLOR;    //显示字符 15mhz
                else
                              pixel_data <= BACK_COLOR;    //显示字符区域的背景色
           end
               else 
                             pixel_data <= BACK_COLOR; 
             12'd1:    
                             if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
                                              && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
                                        if(char_k5k[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
                                           pixel_data <= CHAR_COLOR;    //显示字符 160
                             else
                                           pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                        end
                             else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
                                && (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
                                        if(char_kong10[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
                                           pixel_data <= CHAR_COLOR;    //显示字符 320
                             else
                                           pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                        end
                             else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
                                && (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
                                        if(char_15MHZ[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
                                           pixel_data <= CHAR_COLOR;    //显示字符 15mhz
                             else
                                           pixel_data <= BACK_COLOR;    //显示字符区域的背景色
                        end
                            else 
                                          pixel_data <= BACK_COLOR;  
            default:  if((pixel_xpos >= CHAR_X_START_20 - 1'b1) && (pixel_xpos < CHAR_X_START_20 + CHAR_WIDTH_20 - 1'b1)
            && (pixel_ypos >= CHAR_Y_START_20) && (pixel_ypos < CHAR_Y_START_20 + CHAR_HEIGHT)) begin
      if(char_kong20[y_cnt_20][CHAR_WIDTH_20 -1'b1 - x_cnt_20])
         pixel_data <= CHAR_COLOR;    //显示字符 20
else
         pixel_data <= BACK_COLOR;    //显示字符区域的背景色
end
else if((pixel_xpos >= CHAR_X_START_40 - 1'b1) && (pixel_xpos < CHAR_X_START_40 + CHAR_WIDTH_40 - 1'b1)
&& (pixel_ypos >= CHAR_Y_START_40) && (pixel_ypos < CHAR_Y_START_40 + CHAR_HEIGHT)) begin
      if(char_kong40[y_cnt_40][CHAR_WIDTH_40 -1'b1 - x_cnt_40])
         pixel_data <= CHAR_COLOR;    //显示字符 40
else
         pixel_data <= BACK_COLOR;    //显示字符区域的背景色
end
else if((pixel_xpos >= CHAR_X_START_60 - 1'b1) && (pixel_xpos < CHAR_X_START_60 + CHAR_WIDTH_60 - 1'b1)
&& (pixel_ypos >= CHAR_Y_START_60) && (pixel_ypos < CHAR_Y_START_60 + CHAR_HEIGHT)) begin
      if(char_60KHZ[y_cnt_60][CHAR_WIDTH_60 -1'b1 - x_cnt_60])
         pixel_data <= CHAR_COLOR;    //显示字符 60/KHZ
else
         pixel_data <= BACK_COLOR;    //显示字符区域的背景色
end
else 
   pixel_data <= BACK_COLOR; 
     endcase 
   end 
                





endmodule





